--
-- File            :   symbol_mem_pkg.vhd
-- Autor           :   Vlasov D.V.
-- Data            :   2019.06.10
-- Language        :   VHDL
-- Description     :   This symbol memory file for DebugScreenCore
-- Copyright(c)    :   2019 Vlasov D.V.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library dsc;
use dsc.dsc_mem_pkg.all;

package symbol_mem_pkg is

    constant symbol_mem_hex : mem_t(4095 downto 0)(7 downto 0) :=
    (
           0 => 8X"00",
           1 => 8X"00",
           2 => 8X"00",
           3 => 8X"00",
           4 => 8X"00",
           5 => 8X"00",
           6 => 8X"00",
           7 => 8X"00",
           8 => 8X"00",
           9 => 8X"00",
          10 => 8X"00",
          11 => 8X"00",
          12 => 8X"00",
          13 => 8X"00",
          14 => 8X"00",
          15 => 8X"00",
          16 => 8X"00",
          17 => 8X"00",
          18 => 8X"7E",
          19 => 8X"81",
          20 => 8X"A5",
          21 => 8X"A5",
          22 => 8X"A5",
          23 => 8X"81",
          24 => 8X"81",
          25 => 8X"BD",
          26 => 8X"99",
          27 => 8X"81",
          28 => 8X"7E",
          29 => 8X"00",
          30 => 8X"00",
          31 => 8X"00",
          32 => 8X"00",
          33 => 8X"00",
          34 => 8X"7E",
          35 => 8X"FF",
          36 => 8X"DB",
          37 => 8X"DB",
          38 => 8X"DB",
          39 => 8X"FF",
          40 => 8X"FF",
          41 => 8X"C3",
          42 => 8X"E7",
          43 => 8X"FF",
          44 => 8X"7E",
          45 => 8X"00",
          46 => 8X"00",
          47 => 8X"00",
          48 => 8X"00",
          49 => 8X"00",
          50 => 8X"6C",
          51 => 8X"FE",
          52 => 8X"FE",
          53 => 8X"FE",
          54 => 8X"FE",
          55 => 8X"FE",
          56 => 8X"FE",
          57 => 8X"7C",
          58 => 8X"38",
          59 => 8X"10",
          60 => 8X"00",
          61 => 8X"00",
          62 => 8X"00",
          63 => 8X"00",
          64 => 8X"00",
          65 => 8X"00",
          66 => 8X"00",
          67 => 8X"00",
          68 => 8X"10",
          69 => 8X"38",
          70 => 8X"7C",
          71 => 8X"FE",
          72 => 8X"7C",
          73 => 8X"38",
          74 => 8X"10",
          75 => 8X"00",
          76 => 8X"00",
          77 => 8X"00",
          78 => 8X"00",
          79 => 8X"00",
          80 => 8X"00",
          81 => 8X"00",
          82 => 8X"00",
          83 => 8X"18",
          84 => 8X"3C",
          85 => 8X"3C",
          86 => 8X"E7",
          87 => 8X"E7",
          88 => 8X"E7",
          89 => 8X"18",
          90 => 8X"18",
          91 => 8X"3C",
          92 => 8X"00",
          93 => 8X"00",
          94 => 8X"00",
          95 => 8X"00",
          96 => 8X"00",
          97 => 8X"00",
          98 => 8X"00",
          99 => 8X"18",
         100 => 8X"3C",
         101 => 8X"7E",
         102 => 8X"FF",
         103 => 8X"FF",
         104 => 8X"7E",
         105 => 8X"18",
         106 => 8X"18",
         107 => 8X"3C",
         108 => 8X"00",
         109 => 8X"00",
         110 => 8X"00",
         111 => 8X"00",
         112 => 8X"00",
         113 => 8X"00",
         114 => 8X"00",
         115 => 8X"00",
         116 => 8X"00",
         117 => 8X"18",
         118 => 8X"3C",
         119 => 8X"3C",
         120 => 8X"18",
         121 => 8X"00",
         122 => 8X"00",
         123 => 8X"00",
         124 => 8X"00",
         125 => 8X"00",
         126 => 8X"00",
         127 => 8X"00",
         128 => 8X"FF",
         129 => 8X"FF",
         130 => 8X"FF",
         131 => 8X"FF",
         132 => 8X"FF",
         133 => 8X"FF",
         134 => 8X"E7",
         135 => 8X"C3",
         136 => 8X"C3",
         137 => 8X"E7",
         138 => 8X"FF",
         139 => 8X"FF",
         140 => 8X"FF",
         141 => 8X"FF",
         142 => 8X"FF",
         143 => 8X"FF",
         144 => 8X"00",
         145 => 8X"00",
         146 => 8X"00",
         147 => 8X"00",
         148 => 8X"00",
         149 => 8X"3C",
         150 => 8X"66",
         151 => 8X"42",
         152 => 8X"42",
         153 => 8X"66",
         154 => 8X"3C",
         155 => 8X"00",
         156 => 8X"00",
         157 => 8X"00",
         158 => 8X"00",
         159 => 8X"00",
         160 => 8X"FF",
         161 => 8X"FF",
         162 => 8X"FF",
         163 => 8X"FF",
         164 => 8X"C3",
         165 => 8X"99",
         166 => 8X"BD",
         167 => 8X"BD",
         168 => 8X"99",
         169 => 8X"C3",
         170 => 8X"FF",
         171 => 8X"FF",
         172 => 8X"FF",
         173 => 8X"FF",
         174 => 8X"FF",
         175 => 8X"FF",
         176 => 8X"00",
         177 => 8X"00",
         178 => 8X"00",
         179 => 8X"1E",
         180 => 8X"0E",
         181 => 8X"1A",
         182 => 8X"32",
         183 => 8X"78",
         184 => 8X"CC",
         185 => 8X"CC",
         186 => 8X"CC",
         187 => 8X"78",
         188 => 8X"00",
         189 => 8X"00",
         190 => 8X"00",
         191 => 8X"00",
         192 => 8X"00",
         193 => 8X"00",
         194 => 8X"00",
         195 => 8X"3C",
         196 => 8X"66",
         197 => 8X"66",
         198 => 8X"66",
         199 => 8X"3C",
         200 => 8X"18",
         201 => 8X"7E",
         202 => 8X"18",
         203 => 8X"18",
         204 => 8X"00",
         205 => 8X"00",
         206 => 8X"00",
         207 => 8X"00",
         208 => 8X"00",
         209 => 8X"00",
         210 => 8X"00",
         211 => 8X"3F",
         212 => 8X"33",
         213 => 8X"3F",
         214 => 8X"30",
         215 => 8X"30",
         216 => 8X"30",
         217 => 8X"70",
         218 => 8X"F0",
         219 => 8X"E0",
         220 => 8X"00",
         221 => 8X"00",
         222 => 8X"00",
         223 => 8X"00",
         224 => 8X"00",
         225 => 8X"00",
         226 => 8X"00",
         227 => 8X"7F",
         228 => 8X"63",
         229 => 8X"7F",
         230 => 8X"63",
         231 => 8X"63",
         232 => 8X"63",
         233 => 8X"67",
         234 => 8X"E7",
         235 => 8X"E6",
         236 => 8X"C0",
         237 => 8X"00",
         238 => 8X"00",
         239 => 8X"00",
         240 => 8X"00",
         241 => 8X"00",
         242 => 8X"00",
         243 => 8X"18",
         244 => 8X"18",
         245 => 8X"DB",
         246 => 8X"3C",
         247 => 8X"E7",
         248 => 8X"3C",
         249 => 8X"DB",
         250 => 8X"18",
         251 => 8X"18",
         252 => 8X"00",
         253 => 8X"00",
         254 => 8X"00",
         255 => 8X"00",
         256 => 8X"00",
         257 => 8X"00",
         258 => 8X"00",
         259 => 8X"80",
         260 => 8X"C0",
         261 => 8X"E0",
         262 => 8X"F8",
         263 => 8X"FE",
         264 => 8X"F8",
         265 => 8X"E0",
         266 => 8X"C0",
         267 => 8X"80",
         268 => 8X"00",
         269 => 8X"00",
         270 => 8X"00",
         271 => 8X"00",
         272 => 8X"00",
         273 => 8X"00",
         274 => 8X"00",
         275 => 8X"02",
         276 => 8X"06",
         277 => 8X"0E",
         278 => 8X"3E",
         279 => 8X"FE",
         280 => 8X"3E",
         281 => 8X"0E",
         282 => 8X"06",
         283 => 8X"02",
         284 => 8X"00",
         285 => 8X"00",
         286 => 8X"00",
         287 => 8X"00",
         288 => 8X"00",
         289 => 8X"00",
         290 => 8X"00",
         291 => 8X"18",
         292 => 8X"3C",
         293 => 8X"7E",
         294 => 8X"18",
         295 => 8X"18",
         296 => 8X"18",
         297 => 8X"18",
         298 => 8X"18",
         299 => 8X"18",
         300 => 8X"7E",
         301 => 8X"3C",
         302 => 8X"18",
         303 => 8X"00",
         304 => 8X"00",
         305 => 8X"00",
         306 => 8X"00",
         307 => 8X"66",
         308 => 8X"66",
         309 => 8X"66",
         310 => 8X"66",
         311 => 8X"66",
         312 => 8X"66",
         313 => 8X"00",
         314 => 8X"66",
         315 => 8X"66",
         316 => 8X"00",
         317 => 8X"00",
         318 => 8X"00",
         319 => 8X"00",
         320 => 8X"00",
         321 => 8X"00",
         322 => 8X"00",
         323 => 8X"7F",
         324 => 8X"DB",
         325 => 8X"DB",
         326 => 8X"DB",
         327 => 8X"7B",
         328 => 8X"1B",
         329 => 8X"1B",
         330 => 8X"1B",
         331 => 8X"1B",
         332 => 8X"00",
         333 => 8X"00",
         334 => 8X"00",
         335 => 8X"00",
         336 => 8X"00",
         337 => 8X"00",
         338 => 8X"7C",
         339 => 8X"C6",
         340 => 8X"60",
         341 => 8X"38",
         342 => 8X"6C",
         343 => 8X"C6",
         344 => 8X"C6",
         345 => 8X"6C",
         346 => 8X"38",
         347 => 8X"0C",
         348 => 8X"C6",
         349 => 8X"7C",
         350 => 8X"00",
         351 => 8X"00",
         352 => 8X"00",
         353 => 8X"00",
         354 => 8X"00",
         355 => 8X"00",
         356 => 8X"00",
         357 => 8X"00",
         358 => 8X"00",
         359 => 8X"00",
         360 => 8X"00",
         361 => 8X"FE",
         362 => 8X"FE",
         363 => 8X"FE",
         364 => 8X"00",
         365 => 8X"00",
         366 => 8X"00",
         367 => 8X"00",
         368 => 8X"00",
         369 => 8X"00",
         370 => 8X"00",
         371 => 8X"18",
         372 => 8X"3C",
         373 => 8X"7E",
         374 => 8X"18",
         375 => 8X"18",
         376 => 8X"18",
         377 => 8X"7E",
         378 => 8X"3C",
         379 => 8X"18",
         380 => 8X"7E",
         381 => 8X"00",
         382 => 8X"00",
         383 => 8X"00",
         384 => 8X"00",
         385 => 8X"00",
         386 => 8X"00",
         387 => 8X"18",
         388 => 8X"3C",
         389 => 8X"7E",
         390 => 8X"18",
         391 => 8X"18",
         392 => 8X"18",
         393 => 8X"18",
         394 => 8X"18",
         395 => 8X"18",
         396 => 8X"18",
         397 => 8X"18",
         398 => 8X"18",
         399 => 8X"00",
         400 => 8X"00",
         401 => 8X"00",
         402 => 8X"00",
         403 => 8X"18",
         404 => 8X"18",
         405 => 8X"18",
         406 => 8X"18",
         407 => 8X"18",
         408 => 8X"18",
         409 => 8X"18",
         410 => 8X"18",
         411 => 8X"18",
         412 => 8X"7E",
         413 => 8X"3C",
         414 => 8X"18",
         415 => 8X"00",
         416 => 8X"00",
         417 => 8X"00",
         418 => 8X"00",
         419 => 8X"00",
         420 => 8X"00",
         421 => 8X"18",
         422 => 8X"0C",
         423 => 8X"FE",
         424 => 8X"0C",
         425 => 8X"18",
         426 => 8X"00",
         427 => 8X"00",
         428 => 8X"00",
         429 => 8X"00",
         430 => 8X"00",
         431 => 8X"00",
         432 => 8X"00",
         433 => 8X"00",
         434 => 8X"00",
         435 => 8X"00",
         436 => 8X"00",
         437 => 8X"30",
         438 => 8X"60",
         439 => 8X"FE",
         440 => 8X"60",
         441 => 8X"30",
         442 => 8X"00",
         443 => 8X"00",
         444 => 8X"00",
         445 => 8X"00",
         446 => 8X"00",
         447 => 8X"00",
         448 => 8X"00",
         449 => 8X"00",
         450 => 8X"00",
         451 => 8X"00",
         452 => 8X"00",
         453 => 8X"00",
         454 => 8X"C0",
         455 => 8X"C0",
         456 => 8X"C0",
         457 => 8X"FE",
         458 => 8X"00",
         459 => 8X"00",
         460 => 8X"00",
         461 => 8X"00",
         462 => 8X"00",
         463 => 8X"00",
         464 => 8X"00",
         465 => 8X"00",
         466 => 8X"00",
         467 => 8X"00",
         468 => 8X"00",
         469 => 8X"28",
         470 => 8X"6C",
         471 => 8X"FE",
         472 => 8X"6C",
         473 => 8X"28",
         474 => 8X"00",
         475 => 8X"00",
         476 => 8X"00",
         477 => 8X"00",
         478 => 8X"00",
         479 => 8X"00",
         480 => 8X"00",
         481 => 8X"00",
         482 => 8X"00",
         483 => 8X"00",
         484 => 8X"10",
         485 => 8X"38",
         486 => 8X"38",
         487 => 8X"7C",
         488 => 8X"7C",
         489 => 8X"FE",
         490 => 8X"FE",
         491 => 8X"00",
         492 => 8X"00",
         493 => 8X"00",
         494 => 8X"00",
         495 => 8X"00",
         496 => 8X"00",
         497 => 8X"00",
         498 => 8X"00",
         499 => 8X"FE",
         500 => 8X"7C",
         501 => 8X"38",
         502 => 8X"10",
         503 => 8X"00",
         504 => 8X"00",
         505 => 8X"00",
         506 => 8X"00",
         507 => 8X"00",
         508 => 8X"00",
         509 => 8X"00",
         510 => 8X"00",
         511 => 8X"00",
         512 => 8X"00",
         513 => 8X"00",
         514 => 8X"00",
         515 => 8X"00",
         516 => 8X"00",
         517 => 8X"00",
         518 => 8X"00",
         519 => 8X"00",
         520 => 8X"00",
         521 => 8X"00",
         522 => 8X"00",
         523 => 8X"00",
         524 => 8X"00",
         525 => 8X"00",
         526 => 8X"00",
         527 => 8X"00",
         528 => 8X"00",
         529 => 8X"00",
         530 => 8X"18",
         531 => 8X"3C",
         532 => 8X"3C",
         533 => 8X"3C",
         534 => 8X"3C",
         535 => 8X"18",
         536 => 8X"18",
         537 => 8X"18",
         538 => 8X"00",
         539 => 8X"00",
         540 => 8X"18",
         541 => 8X"00",
         542 => 8X"00",
         543 => 8X"00",
         544 => 8X"00",
         545 => 8X"66",
         546 => 8X"66",
         547 => 8X"66",
         548 => 8X"66",
         549 => 8X"66",
         550 => 8X"24",
         551 => 8X"00",
         552 => 8X"00",
         553 => 8X"00",
         554 => 8X"00",
         555 => 8X"00",
         556 => 8X"00",
         557 => 8X"00",
         558 => 8X"00",
         559 => 8X"00",
         560 => 8X"00",
         561 => 8X"00",
         562 => 8X"6C",
         563 => 8X"6C",
         564 => 8X"6C",
         565 => 8X"FE",
         566 => 8X"6C",
         567 => 8X"6C",
         568 => 8X"6C",
         569 => 8X"FE",
         570 => 8X"6C",
         571 => 8X"6C",
         572 => 8X"6C",
         573 => 8X"00",
         574 => 8X"00",
         575 => 8X"00",
         576 => 8X"18",
         577 => 8X"18",
         578 => 8X"18",
         579 => 8X"7C",
         580 => 8X"C6",
         581 => 8X"C2",
         582 => 8X"C0",
         583 => 8X"7C",
         584 => 8X"06",
         585 => 8X"86",
         586 => 8X"C6",
         587 => 8X"7C",
         588 => 8X"18",
         589 => 8X"18",
         590 => 8X"18",
         591 => 8X"00",
         592 => 8X"00",
         593 => 8X"00",
         594 => 8X"00",
         595 => 8X"00",
         596 => 8X"00",
         597 => 8X"C2",
         598 => 8X"C6",
         599 => 8X"0C",
         600 => 8X"18",
         601 => 8X"30",
         602 => 8X"66",
         603 => 8X"C6",
         604 => 8X"00",
         605 => 8X"00",
         606 => 8X"00",
         607 => 8X"00",
         608 => 8X"00",
         609 => 8X"00",
         610 => 8X"38",
         611 => 8X"6C",
         612 => 8X"6C",
         613 => 8X"6C",
         614 => 8X"38",
         615 => 8X"76",
         616 => 8X"DC",
         617 => 8X"CC",
         618 => 8X"CC",
         619 => 8X"CC",
         620 => 8X"76",
         621 => 8X"00",
         622 => 8X"00",
         623 => 8X"00",
         624 => 8X"00",
         625 => 8X"30",
         626 => 8X"30",
         627 => 8X"30",
         628 => 8X"30",
         629 => 8X"60",
         630 => 8X"00",
         631 => 8X"00",
         632 => 8X"00",
         633 => 8X"00",
         634 => 8X"00",
         635 => 8X"00",
         636 => 8X"00",
         637 => 8X"00",
         638 => 8X"00",
         639 => 8X"00",
         640 => 8X"00",
         641 => 8X"00",
         642 => 8X"0C",
         643 => 8X"18",
         644 => 8X"30",
         645 => 8X"30",
         646 => 8X"30",
         647 => 8X"30",
         648 => 8X"30",
         649 => 8X"30",
         650 => 8X"30",
         651 => 8X"18",
         652 => 8X"0C",
         653 => 8X"00",
         654 => 8X"00",
         655 => 8X"00",
         656 => 8X"00",
         657 => 8X"00",
         658 => 8X"30",
         659 => 8X"18",
         660 => 8X"0C",
         661 => 8X"0C",
         662 => 8X"0C",
         663 => 8X"0C",
         664 => 8X"0C",
         665 => 8X"0C",
         666 => 8X"0C",
         667 => 8X"18",
         668 => 8X"30",
         669 => 8X"00",
         670 => 8X"00",
         671 => 8X"00",
         672 => 8X"00",
         673 => 8X"00",
         674 => 8X"00",
         675 => 8X"00",
         676 => 8X"66",
         677 => 8X"66",
         678 => 8X"3C",
         679 => 8X"FF",
         680 => 8X"3C",
         681 => 8X"66",
         682 => 8X"66",
         683 => 8X"00",
         684 => 8X"00",
         685 => 8X"00",
         686 => 8X"00",
         687 => 8X"00",
         688 => 8X"00",
         689 => 8X"00",
         690 => 8X"00",
         691 => 8X"00",
         692 => 8X"18",
         693 => 8X"18",
         694 => 8X"18",
         695 => 8X"7E",
         696 => 8X"18",
         697 => 8X"18",
         698 => 8X"18",
         699 => 8X"00",
         700 => 8X"00",
         701 => 8X"00",
         702 => 8X"00",
         703 => 8X"00",
         704 => 8X"00",
         705 => 8X"00",
         706 => 8X"00",
         707 => 8X"00",
         708 => 8X"00",
         709 => 8X"00",
         710 => 8X"00",
         711 => 8X"00",
         712 => 8X"00",
         713 => 8X"18",
         714 => 8X"18",
         715 => 8X"18",
         716 => 8X"18",
         717 => 8X"30",
         718 => 8X"00",
         719 => 8X"00",
         720 => 8X"00",
         721 => 8X"00",
         722 => 8X"00",
         723 => 8X"00",
         724 => 8X"00",
         725 => 8X"00",
         726 => 8X"00",
         727 => 8X"FE",
         728 => 8X"00",
         729 => 8X"00",
         730 => 8X"00",
         731 => 8X"00",
         732 => 8X"00",
         733 => 8X"00",
         734 => 8X"00",
         735 => 8X"00",
         736 => 8X"00",
         737 => 8X"00",
         738 => 8X"00",
         739 => 8X"00",
         740 => 8X"00",
         741 => 8X"00",
         742 => 8X"00",
         743 => 8X"00",
         744 => 8X"00",
         745 => 8X"00",
         746 => 8X"00",
         747 => 8X"18",
         748 => 8X"18",
         749 => 8X"00",
         750 => 8X"00",
         751 => 8X"00",
         752 => 8X"00",
         753 => 8X"00",
         754 => 8X"00",
         755 => 8X"02",
         756 => 8X"06",
         757 => 8X"0C",
         758 => 8X"18",
         759 => 8X"30",
         760 => 8X"60",
         761 => 8X"C0",
         762 => 8X"80",
         763 => 8X"00",
         764 => 8X"00",
         765 => 8X"00",
         766 => 8X"00",
         767 => 8X"00",
         768 => 8X"00",
         769 => 8X"00",
         770 => 8X"7C",
         771 => 8X"C6",
         772 => 8X"C6",
         773 => 8X"CE",
         774 => 8X"DE",
         775 => 8X"F6",
         776 => 8X"F6",
         777 => 8X"E6",
         778 => 8X"C6",
         779 => 8X"C6",
         780 => 8X"7C",
         781 => 8X"00",
         782 => 8X"00",
         783 => 8X"00",
         784 => 8X"00",
         785 => 8X"00",
         786 => 8X"18",
         787 => 8X"18",
         788 => 8X"38",
         789 => 8X"78",
         790 => 8X"18",
         791 => 8X"18",
         792 => 8X"18",
         793 => 8X"18",
         794 => 8X"18",
         795 => 8X"18",
         796 => 8X"7E",
         797 => 8X"00",
         798 => 8X"00",
         799 => 8X"00",
         800 => 8X"00",
         801 => 8X"00",
         802 => 8X"7C",
         803 => 8X"C6",
         804 => 8X"C6",
         805 => 8X"06",
         806 => 8X"06",
         807 => 8X"0C",
         808 => 8X"18",
         809 => 8X"30",
         810 => 8X"60",
         811 => 8X"C6",
         812 => 8X"FE",
         813 => 8X"00",
         814 => 8X"00",
         815 => 8X"00",
         816 => 8X"00",
         817 => 8X"00",
         818 => 8X"7C",
         819 => 8X"C6",
         820 => 8X"06",
         821 => 8X"06",
         822 => 8X"06",
         823 => 8X"3C",
         824 => 8X"06",
         825 => 8X"06",
         826 => 8X"06",
         827 => 8X"C6",
         828 => 8X"7C",
         829 => 8X"00",
         830 => 8X"00",
         831 => 8X"00",
         832 => 8X"00",
         833 => 8X"00",
         834 => 8X"0C",
         835 => 8X"1C",
         836 => 8X"3C",
         837 => 8X"6C",
         838 => 8X"CC",
         839 => 8X"CC",
         840 => 8X"FE",
         841 => 8X"0C",
         842 => 8X"0C",
         843 => 8X"0C",
         844 => 8X"1E",
         845 => 8X"00",
         846 => 8X"00",
         847 => 8X"00",
         848 => 8X"00",
         849 => 8X"00",
         850 => 8X"FE",
         851 => 8X"C0",
         852 => 8X"C0",
         853 => 8X"C0",
         854 => 8X"FC",
         855 => 8X"06",
         856 => 8X"06",
         857 => 8X"06",
         858 => 8X"06",
         859 => 8X"C6",
         860 => 8X"7C",
         861 => 8X"00",
         862 => 8X"00",
         863 => 8X"00",
         864 => 8X"00",
         865 => 8X"00",
         866 => 8X"38",
         867 => 8X"60",
         868 => 8X"C0",
         869 => 8X"C0",
         870 => 8X"FC",
         871 => 8X"C6",
         872 => 8X"C6",
         873 => 8X"C6",
         874 => 8X"C6",
         875 => 8X"C6",
         876 => 8X"7C",
         877 => 8X"00",
         878 => 8X"00",
         879 => 8X"00",
         880 => 8X"00",
         881 => 8X"00",
         882 => 8X"FE",
         883 => 8X"C6",
         884 => 8X"C6",
         885 => 8X"06",
         886 => 8X"06",
         887 => 8X"0C",
         888 => 8X"18",
         889 => 8X"30",
         890 => 8X"30",
         891 => 8X"30",
         892 => 8X"30",
         893 => 8X"00",
         894 => 8X"00",
         895 => 8X"00",
         896 => 8X"00",
         897 => 8X"00",
         898 => 8X"7C",
         899 => 8X"C6",
         900 => 8X"C6",
         901 => 8X"C6",
         902 => 8X"C6",
         903 => 8X"7C",
         904 => 8X"C6",
         905 => 8X"C6",
         906 => 8X"C6",
         907 => 8X"C6",
         908 => 8X"7C",
         909 => 8X"00",
         910 => 8X"00",
         911 => 8X"00",
         912 => 8X"00",
         913 => 8X"00",
         914 => 8X"7C",
         915 => 8X"C6",
         916 => 8X"C6",
         917 => 8X"C6",
         918 => 8X"C6",
         919 => 8X"C6",
         920 => 8X"7E",
         921 => 8X"06",
         922 => 8X"06",
         923 => 8X"0C",
         924 => 8X"78",
         925 => 8X"00",
         926 => 8X"00",
         927 => 8X"00",
         928 => 8X"00",
         929 => 8X"00",
         930 => 8X"00",
         931 => 8X"18",
         932 => 8X"18",
         933 => 8X"00",
         934 => 8X"00",
         935 => 8X"00",
         936 => 8X"00",
         937 => 8X"00",
         938 => 8X"00",
         939 => 8X"18",
         940 => 8X"18",
         941 => 8X"00",
         942 => 8X"00",
         943 => 8X"00",
         944 => 8X"00",
         945 => 8X"00",
         946 => 8X"00",
         947 => 8X"18",
         948 => 8X"18",
         949 => 8X"00",
         950 => 8X"00",
         951 => 8X"00",
         952 => 8X"00",
         953 => 8X"18",
         954 => 8X"18",
         955 => 8X"18",
         956 => 8X"18",
         957 => 8X"30",
         958 => 8X"00",
         959 => 8X"00",
         960 => 8X"00",
         961 => 8X"00",
         962 => 8X"00",
         963 => 8X"06",
         964 => 8X"0C",
         965 => 8X"18",
         966 => 8X"30",
         967 => 8X"60",
         968 => 8X"30",
         969 => 8X"18",
         970 => 8X"0C",
         971 => 8X"06",
         972 => 8X"00",
         973 => 8X"00",
         974 => 8X"00",
         975 => 8X"00",
         976 => 8X"00",
         977 => 8X"00",
         978 => 8X"00",
         979 => 8X"00",
         980 => 8X"00",
         981 => 8X"00",
         982 => 8X"7E",
         983 => 8X"00",
         984 => 8X"00",
         985 => 8X"7E",
         986 => 8X"00",
         987 => 8X"00",
         988 => 8X"00",
         989 => 8X"00",
         990 => 8X"00",
         991 => 8X"00",
         992 => 8X"00",
         993 => 8X"00",
         994 => 8X"00",
         995 => 8X"60",
         996 => 8X"30",
         997 => 8X"18",
         998 => 8X"0C",
         999 => 8X"06",
        1000 => 8X"0C",
        1001 => 8X"18",
        1002 => 8X"30",
        1003 => 8X"60",
        1004 => 8X"00",
        1005 => 8X"00",
        1006 => 8X"00",
        1007 => 8X"00",
        1008 => 8X"00",
        1009 => 8X"00",
        1010 => 8X"7C",
        1011 => 8X"C6",
        1012 => 8X"C6",
        1013 => 8X"C6",
        1014 => 8X"0C",
        1015 => 8X"18",
        1016 => 8X"18",
        1017 => 8X"18",
        1018 => 8X"00",
        1019 => 8X"18",
        1020 => 8X"18",
        1021 => 8X"00",
        1022 => 8X"00",
        1023 => 8X"00",
        1024 => 8X"00",
        1025 => 8X"00",
        1026 => 8X"7C",
        1027 => 8X"C6",
        1028 => 8X"C6",
        1029 => 8X"C6",
        1030 => 8X"DE",
        1031 => 8X"DE",
        1032 => 8X"DE",
        1033 => 8X"DC",
        1034 => 8X"C0",
        1035 => 8X"C0",
        1036 => 8X"7C",
        1037 => 8X"00",
        1038 => 8X"00",
        1039 => 8X"00",
        1040 => 8X"00",
        1041 => 8X"00",
        1042 => 8X"10",
        1043 => 8X"38",
        1044 => 8X"6C",
        1045 => 8X"C6",
        1046 => 8X"C6",
        1047 => 8X"C6",
        1048 => 8X"FE",
        1049 => 8X"C6",
        1050 => 8X"C6",
        1051 => 8X"C6",
        1052 => 8X"C6",
        1053 => 8X"00",
        1054 => 8X"00",
        1055 => 8X"00",
        1056 => 8X"00",
        1057 => 8X"00",
        1058 => 8X"FC",
        1059 => 8X"66",
        1060 => 8X"66",
        1061 => 8X"66",
        1062 => 8X"66",
        1063 => 8X"7C",
        1064 => 8X"66",
        1065 => 8X"66",
        1066 => 8X"66",
        1067 => 8X"66",
        1068 => 8X"FC",
        1069 => 8X"00",
        1070 => 8X"00",
        1071 => 8X"00",
        1072 => 8X"00",
        1073 => 8X"00",
        1074 => 8X"7C",
        1075 => 8X"C6",
        1076 => 8X"C6",
        1077 => 8X"C0",
        1078 => 8X"C0",
        1079 => 8X"C0",
        1080 => 8X"C0",
        1081 => 8X"C6",
        1082 => 8X"C6",
        1083 => 8X"C6",
        1084 => 8X"7C",
        1085 => 8X"00",
        1086 => 8X"00",
        1087 => 8X"00",
        1088 => 8X"00",
        1089 => 8X"00",
        1090 => 8X"FC",
        1091 => 8X"66",
        1092 => 8X"66",
        1093 => 8X"66",
        1094 => 8X"66",
        1095 => 8X"66",
        1096 => 8X"66",
        1097 => 8X"66",
        1098 => 8X"66",
        1099 => 8X"66",
        1100 => 8X"FC",
        1101 => 8X"00",
        1102 => 8X"00",
        1103 => 8X"00",
        1104 => 8X"00",
        1105 => 8X"00",
        1106 => 8X"FE",
        1107 => 8X"66",
        1108 => 8X"62",
        1109 => 8X"60",
        1110 => 8X"68",
        1111 => 8X"78",
        1112 => 8X"68",
        1113 => 8X"68",
        1114 => 8X"62",
        1115 => 8X"66",
        1116 => 8X"FE",
        1117 => 8X"00",
        1118 => 8X"00",
        1119 => 8X"00",
        1120 => 8X"00",
        1121 => 8X"00",
        1122 => 8X"FE",
        1123 => 8X"66",
        1124 => 8X"62",
        1125 => 8X"60",
        1126 => 8X"68",
        1127 => 8X"78",
        1128 => 8X"68",
        1129 => 8X"68",
        1130 => 8X"60",
        1131 => 8X"60",
        1132 => 8X"F0",
        1133 => 8X"00",
        1134 => 8X"00",
        1135 => 8X"00",
        1136 => 8X"00",
        1137 => 8X"00",
        1138 => 8X"7C",
        1139 => 8X"C6",
        1140 => 8X"C6",
        1141 => 8X"C0",
        1142 => 8X"C0",
        1143 => 8X"C0",
        1144 => 8X"DE",
        1145 => 8X"C6",
        1146 => 8X"C6",
        1147 => 8X"C6",
        1148 => 8X"7C",
        1149 => 8X"00",
        1150 => 8X"00",
        1151 => 8X"00",
        1152 => 8X"00",
        1153 => 8X"00",
        1154 => 8X"C6",
        1155 => 8X"C6",
        1156 => 8X"C6",
        1157 => 8X"C6",
        1158 => 8X"C6",
        1159 => 8X"FE",
        1160 => 8X"C6",
        1161 => 8X"C6",
        1162 => 8X"C6",
        1163 => 8X"C6",
        1164 => 8X"C6",
        1165 => 8X"00",
        1166 => 8X"00",
        1167 => 8X"00",
        1168 => 8X"00",
        1169 => 8X"00",
        1170 => 8X"3C",
        1171 => 8X"18",
        1172 => 8X"18",
        1173 => 8X"18",
        1174 => 8X"18",
        1175 => 8X"18",
        1176 => 8X"18",
        1177 => 8X"18",
        1178 => 8X"18",
        1179 => 8X"18",
        1180 => 8X"3C",
        1181 => 8X"00",
        1182 => 8X"00",
        1183 => 8X"00",
        1184 => 8X"00",
        1185 => 8X"00",
        1186 => 8X"1E",
        1187 => 8X"0C",
        1188 => 8X"0C",
        1189 => 8X"0C",
        1190 => 8X"0C",
        1191 => 8X"0C",
        1192 => 8X"0C",
        1193 => 8X"0C",
        1194 => 8X"CC",
        1195 => 8X"CC",
        1196 => 8X"78",
        1197 => 8X"00",
        1198 => 8X"00",
        1199 => 8X"00",
        1200 => 8X"00",
        1201 => 8X"00",
        1202 => 8X"E6",
        1203 => 8X"66",
        1204 => 8X"66",
        1205 => 8X"6C",
        1206 => 8X"6C",
        1207 => 8X"78",
        1208 => 8X"6C",
        1209 => 8X"6C",
        1210 => 8X"66",
        1211 => 8X"66",
        1212 => 8X"E6",
        1213 => 8X"00",
        1214 => 8X"00",
        1215 => 8X"00",
        1216 => 8X"00",
        1217 => 8X"00",
        1218 => 8X"F0",
        1219 => 8X"60",
        1220 => 8X"60",
        1221 => 8X"60",
        1222 => 8X"60",
        1223 => 8X"60",
        1224 => 8X"60",
        1225 => 8X"60",
        1226 => 8X"62",
        1227 => 8X"66",
        1228 => 8X"FE",
        1229 => 8X"00",
        1230 => 8X"00",
        1231 => 8X"00",
        1232 => 8X"00",
        1233 => 8X"00",
        1234 => 8X"C6",
        1235 => 8X"C6",
        1236 => 8X"EE",
        1237 => 8X"FE",
        1238 => 8X"FE",
        1239 => 8X"D6",
        1240 => 8X"C6",
        1241 => 8X"C6",
        1242 => 8X"C6",
        1243 => 8X"C6",
        1244 => 8X"C6",
        1245 => 8X"00",
        1246 => 8X"00",
        1247 => 8X"00",
        1248 => 8X"00",
        1249 => 8X"00",
        1250 => 8X"C6",
        1251 => 8X"C6",
        1252 => 8X"E6",
        1253 => 8X"F6",
        1254 => 8X"FE",
        1255 => 8X"DE",
        1256 => 8X"CE",
        1257 => 8X"C6",
        1258 => 8X"C6",
        1259 => 8X"C6",
        1260 => 8X"C6",
        1261 => 8X"00",
        1262 => 8X"00",
        1263 => 8X"00",
        1264 => 8X"00",
        1265 => 8X"00",
        1266 => 8X"7C",
        1267 => 8X"C6",
        1268 => 8X"C6",
        1269 => 8X"C6",
        1270 => 8X"C6",
        1271 => 8X"C6",
        1272 => 8X"C6",
        1273 => 8X"C6",
        1274 => 8X"C6",
        1275 => 8X"C6",
        1276 => 8X"7C",
        1277 => 8X"00",
        1278 => 8X"00",
        1279 => 8X"00",
        1280 => 8X"00",
        1281 => 8X"00",
        1282 => 8X"FC",
        1283 => 8X"66",
        1284 => 8X"66",
        1285 => 8X"66",
        1286 => 8X"66",
        1287 => 8X"66",
        1288 => 8X"7C",
        1289 => 8X"60",
        1290 => 8X"60",
        1291 => 8X"60",
        1292 => 8X"F0",
        1293 => 8X"00",
        1294 => 8X"00",
        1295 => 8X"00",
        1296 => 8X"00",
        1297 => 8X"00",
        1298 => 8X"7C",
        1299 => 8X"C6",
        1300 => 8X"C6",
        1301 => 8X"C6",
        1302 => 8X"C6",
        1303 => 8X"C6",
        1304 => 8X"C6",
        1305 => 8X"D6",
        1306 => 8X"DE",
        1307 => 8X"7C",
        1308 => 8X"0C",
        1309 => 8X"00",
        1310 => 8X"00",
        1311 => 8X"00",
        1312 => 8X"00",
        1313 => 8X"00",
        1314 => 8X"FC",
        1315 => 8X"66",
        1316 => 8X"66",
        1317 => 8X"66",
        1318 => 8X"66",
        1319 => 8X"7C",
        1320 => 8X"6C",
        1321 => 8X"66",
        1322 => 8X"66",
        1323 => 8X"66",
        1324 => 8X"E6",
        1325 => 8X"00",
        1326 => 8X"00",
        1327 => 8X"00",
        1328 => 8X"00",
        1329 => 8X"00",
        1330 => 8X"7C",
        1331 => 8X"C6",
        1332 => 8X"C6",
        1333 => 8X"C6",
        1334 => 8X"60",
        1335 => 8X"38",
        1336 => 8X"0C",
        1337 => 8X"C6",
        1338 => 8X"C6",
        1339 => 8X"C6",
        1340 => 8X"7C",
        1341 => 8X"00",
        1342 => 8X"00",
        1343 => 8X"00",
        1344 => 8X"00",
        1345 => 8X"00",
        1346 => 8X"7E",
        1347 => 8X"7E",
        1348 => 8X"5A",
        1349 => 8X"18",
        1350 => 8X"18",
        1351 => 8X"18",
        1352 => 8X"18",
        1353 => 8X"18",
        1354 => 8X"18",
        1355 => 8X"18",
        1356 => 8X"3C",
        1357 => 8X"00",
        1358 => 8X"00",
        1359 => 8X"00",
        1360 => 8X"00",
        1361 => 8X"00",
        1362 => 8X"C6",
        1363 => 8X"C6",
        1364 => 8X"C6",
        1365 => 8X"C6",
        1366 => 8X"C6",
        1367 => 8X"C6",
        1368 => 8X"C6",
        1369 => 8X"C6",
        1370 => 8X"C6",
        1371 => 8X"C6",
        1372 => 8X"7C",
        1373 => 8X"00",
        1374 => 8X"00",
        1375 => 8X"00",
        1376 => 8X"00",
        1377 => 8X"00",
        1378 => 8X"C6",
        1379 => 8X"C6",
        1380 => 8X"C6",
        1381 => 8X"C6",
        1382 => 8X"C6",
        1383 => 8X"C6",
        1384 => 8X"C6",
        1385 => 8X"C6",
        1386 => 8X"6C",
        1387 => 8X"38",
        1388 => 8X"10",
        1389 => 8X"00",
        1390 => 8X"00",
        1391 => 8X"00",
        1392 => 8X"00",
        1393 => 8X"00",
        1394 => 8X"C6",
        1395 => 8X"C6",
        1396 => 8X"C6",
        1397 => 8X"C6",
        1398 => 8X"C6",
        1399 => 8X"D6",
        1400 => 8X"D6",
        1401 => 8X"FE",
        1402 => 8X"7C",
        1403 => 8X"6C",
        1404 => 8X"6C",
        1405 => 8X"00",
        1406 => 8X"00",
        1407 => 8X"00",
        1408 => 8X"00",
        1409 => 8X"00",
        1410 => 8X"C6",
        1411 => 8X"C6",
        1412 => 8X"C6",
        1413 => 8X"6C",
        1414 => 8X"38",
        1415 => 8X"38",
        1416 => 8X"38",
        1417 => 8X"6C",
        1418 => 8X"C6",
        1419 => 8X"C6",
        1420 => 8X"C6",
        1421 => 8X"00",
        1422 => 8X"00",
        1423 => 8X"00",
        1424 => 8X"00",
        1425 => 8X"00",
        1426 => 8X"66",
        1427 => 8X"66",
        1428 => 8X"66",
        1429 => 8X"66",
        1430 => 8X"66",
        1431 => 8X"3C",
        1432 => 8X"18",
        1433 => 8X"18",
        1434 => 8X"18",
        1435 => 8X"18",
        1436 => 8X"3C",
        1437 => 8X"00",
        1438 => 8X"00",
        1439 => 8X"00",
        1440 => 8X"00",
        1441 => 8X"00",
        1442 => 8X"FE",
        1443 => 8X"C6",
        1444 => 8X"C6",
        1445 => 8X"8C",
        1446 => 8X"18",
        1447 => 8X"30",
        1448 => 8X"60",
        1449 => 8X"C2",
        1450 => 8X"C6",
        1451 => 8X"C6",
        1452 => 8X"FE",
        1453 => 8X"00",
        1454 => 8X"00",
        1455 => 8X"00",
        1456 => 8X"00",
        1457 => 8X"00",
        1458 => 8X"3C",
        1459 => 8X"30",
        1460 => 8X"30",
        1461 => 8X"30",
        1462 => 8X"30",
        1463 => 8X"30",
        1464 => 8X"30",
        1465 => 8X"30",
        1466 => 8X"30",
        1467 => 8X"30",
        1468 => 8X"3C",
        1469 => 8X"00",
        1470 => 8X"00",
        1471 => 8X"00",
        1472 => 8X"00",
        1473 => 8X"00",
        1474 => 8X"00",
        1475 => 8X"80",
        1476 => 8X"C0",
        1477 => 8X"E0",
        1478 => 8X"70",
        1479 => 8X"38",
        1480 => 8X"1C",
        1481 => 8X"0E",
        1482 => 8X"06",
        1483 => 8X"02",
        1484 => 8X"00",
        1485 => 8X"00",
        1486 => 8X"00",
        1487 => 8X"00",
        1488 => 8X"00",
        1489 => 8X"00",
        1490 => 8X"3C",
        1491 => 8X"0C",
        1492 => 8X"0C",
        1493 => 8X"0C",
        1494 => 8X"0C",
        1495 => 8X"0C",
        1496 => 8X"0C",
        1497 => 8X"0C",
        1498 => 8X"0C",
        1499 => 8X"0C",
        1500 => 8X"3C",
        1501 => 8X"00",
        1502 => 8X"00",
        1503 => 8X"00",
        1504 => 8X"10",
        1505 => 8X"10",
        1506 => 8X"38",
        1507 => 8X"6C",
        1508 => 8X"C6",
        1509 => 8X"00",
        1510 => 8X"00",
        1511 => 8X"00",
        1512 => 8X"00",
        1513 => 8X"00",
        1514 => 8X"00",
        1515 => 8X"00",
        1516 => 8X"00",
        1517 => 8X"00",
        1518 => 8X"00",
        1519 => 8X"00",
        1520 => 8X"00",
        1521 => 8X"00",
        1522 => 8X"00",
        1523 => 8X"00",
        1524 => 8X"00",
        1525 => 8X"00",
        1526 => 8X"00",
        1527 => 8X"00",
        1528 => 8X"00",
        1529 => 8X"00",
        1530 => 8X"00",
        1531 => 8X"00",
        1532 => 8X"00",
        1533 => 8X"FF",
        1534 => 8X"FF",
        1535 => 8X"00",
        1536 => 8X"30",
        1537 => 8X"30",
        1538 => 8X"30",
        1539 => 8X"18",
        1540 => 8X"00",
        1541 => 8X"00",
        1542 => 8X"00",
        1543 => 8X"00",
        1544 => 8X"00",
        1545 => 8X"00",
        1546 => 8X"00",
        1547 => 8X"00",
        1548 => 8X"00",
        1549 => 8X"00",
        1550 => 8X"00",
        1551 => 8X"00",
        1552 => 8X"00",
        1553 => 8X"00",
        1554 => 8X"00",
        1555 => 8X"00",
        1556 => 8X"00",
        1557 => 8X"78",
        1558 => 8X"CC",
        1559 => 8X"0C",
        1560 => 8X"7C",
        1561 => 8X"CC",
        1562 => 8X"CC",
        1563 => 8X"CC",
        1564 => 8X"76",
        1565 => 8X"00",
        1566 => 8X"00",
        1567 => 8X"00",
        1568 => 8X"00",
        1569 => 8X"00",
        1570 => 8X"E0",
        1571 => 8X"60",
        1572 => 8X"60",
        1573 => 8X"60",
        1574 => 8X"78",
        1575 => 8X"6C",
        1576 => 8X"66",
        1577 => 8X"66",
        1578 => 8X"66",
        1579 => 8X"66",
        1580 => 8X"7C",
        1581 => 8X"00",
        1582 => 8X"00",
        1583 => 8X"00",
        1584 => 8X"00",
        1585 => 8X"00",
        1586 => 8X"00",
        1587 => 8X"00",
        1588 => 8X"00",
        1589 => 8X"7C",
        1590 => 8X"C6",
        1591 => 8X"C6",
        1592 => 8X"C0",
        1593 => 8X"C0",
        1594 => 8X"C6",
        1595 => 8X"C6",
        1596 => 8X"7C",
        1597 => 8X"00",
        1598 => 8X"00",
        1599 => 8X"00",
        1600 => 8X"00",
        1601 => 8X"00",
        1602 => 8X"1C",
        1603 => 8X"0C",
        1604 => 8X"0C",
        1605 => 8X"0C",
        1606 => 8X"3C",
        1607 => 8X"6C",
        1608 => 8X"CC",
        1609 => 8X"CC",
        1610 => 8X"CC",
        1611 => 8X"CC",
        1612 => 8X"76",
        1613 => 8X"00",
        1614 => 8X"00",
        1615 => 8X"00",
        1616 => 8X"00",
        1617 => 8X"00",
        1618 => 8X"00",
        1619 => 8X"00",
        1620 => 8X"00",
        1621 => 8X"7C",
        1622 => 8X"C6",
        1623 => 8X"C6",
        1624 => 8X"FE",
        1625 => 8X"C0",
        1626 => 8X"C6",
        1627 => 8X"C6",
        1628 => 8X"7C",
        1629 => 8X"00",
        1630 => 8X"00",
        1631 => 8X"00",
        1632 => 8X"00",
        1633 => 8X"00",
        1634 => 8X"38",
        1635 => 8X"6C",
        1636 => 8X"64",
        1637 => 8X"60",
        1638 => 8X"F0",
        1639 => 8X"60",
        1640 => 8X"60",
        1641 => 8X"60",
        1642 => 8X"60",
        1643 => 8X"60",
        1644 => 8X"F0",
        1645 => 8X"00",
        1646 => 8X"00",
        1647 => 8X"00",
        1648 => 8X"00",
        1649 => 8X"00",
        1650 => 8X"00",
        1651 => 8X"00",
        1652 => 8X"00",
        1653 => 8X"76",
        1654 => 8X"CC",
        1655 => 8X"CC",
        1656 => 8X"CC",
        1657 => 8X"CC",
        1658 => 8X"CC",
        1659 => 8X"7C",
        1660 => 8X"0C",
        1661 => 8X"CC",
        1662 => 8X"78",
        1663 => 8X"00",
        1664 => 8X"00",
        1665 => 8X"00",
        1666 => 8X"E0",
        1667 => 8X"60",
        1668 => 8X"60",
        1669 => 8X"6C",
        1670 => 8X"76",
        1671 => 8X"66",
        1672 => 8X"66",
        1673 => 8X"66",
        1674 => 8X"66",
        1675 => 8X"66",
        1676 => 8X"E6",
        1677 => 8X"00",
        1678 => 8X"00",
        1679 => 8X"00",
        1680 => 8X"00",
        1681 => 8X"00",
        1682 => 8X"18",
        1683 => 8X"18",
        1684 => 8X"00",
        1685 => 8X"38",
        1686 => 8X"18",
        1687 => 8X"18",
        1688 => 8X"18",
        1689 => 8X"18",
        1690 => 8X"18",
        1691 => 8X"18",
        1692 => 8X"3C",
        1693 => 8X"00",
        1694 => 8X"00",
        1695 => 8X"00",
        1696 => 8X"00",
        1697 => 8X"00",
        1698 => 8X"06",
        1699 => 8X"06",
        1700 => 8X"00",
        1701 => 8X"0E",
        1702 => 8X"06",
        1703 => 8X"06",
        1704 => 8X"06",
        1705 => 8X"06",
        1706 => 8X"06",
        1707 => 8X"06",
        1708 => 8X"66",
        1709 => 8X"66",
        1710 => 8X"3C",
        1711 => 8X"00",
        1712 => 8X"00",
        1713 => 8X"00",
        1714 => 8X"E0",
        1715 => 8X"60",
        1716 => 8X"60",
        1717 => 8X"66",
        1718 => 8X"66",
        1719 => 8X"6C",
        1720 => 8X"78",
        1721 => 8X"6C",
        1722 => 8X"66",
        1723 => 8X"66",
        1724 => 8X"E6",
        1725 => 8X"00",
        1726 => 8X"00",
        1727 => 8X"00",
        1728 => 8X"00",
        1729 => 8X"00",
        1730 => 8X"38",
        1731 => 8X"18",
        1732 => 8X"18",
        1733 => 8X"18",
        1734 => 8X"18",
        1735 => 8X"18",
        1736 => 8X"18",
        1737 => 8X"18",
        1738 => 8X"18",
        1739 => 8X"18",
        1740 => 8X"3C",
        1741 => 8X"00",
        1742 => 8X"00",
        1743 => 8X"00",
        1744 => 8X"00",
        1745 => 8X"00",
        1746 => 8X"00",
        1747 => 8X"00",
        1748 => 8X"00",
        1749 => 8X"EC",
        1750 => 8X"FE",
        1751 => 8X"D6",
        1752 => 8X"D6",
        1753 => 8X"D6",
        1754 => 8X"C6",
        1755 => 8X"C6",
        1756 => 8X"C6",
        1757 => 8X"00",
        1758 => 8X"00",
        1759 => 8X"00",
        1760 => 8X"00",
        1761 => 8X"00",
        1762 => 8X"00",
        1763 => 8X"00",
        1764 => 8X"00",
        1765 => 8X"DC",
        1766 => 8X"66",
        1767 => 8X"66",
        1768 => 8X"66",
        1769 => 8X"66",
        1770 => 8X"66",
        1771 => 8X"66",
        1772 => 8X"66",
        1773 => 8X"00",
        1774 => 8X"00",
        1775 => 8X"00",
        1776 => 8X"00",
        1777 => 8X"00",
        1778 => 8X"00",
        1779 => 8X"00",
        1780 => 8X"00",
        1781 => 8X"7C",
        1782 => 8X"C6",
        1783 => 8X"C6",
        1784 => 8X"C6",
        1785 => 8X"C6",
        1786 => 8X"C6",
        1787 => 8X"C6",
        1788 => 8X"7C",
        1789 => 8X"00",
        1790 => 8X"00",
        1791 => 8X"00",
        1792 => 8X"00",
        1793 => 8X"00",
        1794 => 8X"00",
        1795 => 8X"00",
        1796 => 8X"00",
        1797 => 8X"DC",
        1798 => 8X"66",
        1799 => 8X"66",
        1800 => 8X"66",
        1801 => 8X"66",
        1802 => 8X"66",
        1803 => 8X"66",
        1804 => 8X"7C",
        1805 => 8X"60",
        1806 => 8X"F0",
        1807 => 8X"00",
        1808 => 8X"00",
        1809 => 8X"00",
        1810 => 8X"00",
        1811 => 8X"00",
        1812 => 8X"00",
        1813 => 8X"76",
        1814 => 8X"CC",
        1815 => 8X"CC",
        1816 => 8X"CC",
        1817 => 8X"CC",
        1818 => 8X"CC",
        1819 => 8X"CC",
        1820 => 8X"7C",
        1821 => 8X"0C",
        1822 => 8X"1E",
        1823 => 8X"00",
        1824 => 8X"00",
        1825 => 8X"00",
        1826 => 8X"00",
        1827 => 8X"00",
        1828 => 8X"00",
        1829 => 8X"DC",
        1830 => 8X"76",
        1831 => 8X"66",
        1832 => 8X"60",
        1833 => 8X"60",
        1834 => 8X"60",
        1835 => 8X"60",
        1836 => 8X"F0",
        1837 => 8X"00",
        1838 => 8X"00",
        1839 => 8X"00",
        1840 => 8X"00",
        1841 => 8X"00",
        1842 => 8X"00",
        1843 => 8X"00",
        1844 => 8X"00",
        1845 => 8X"7C",
        1846 => 8X"C6",
        1847 => 8X"C6",
        1848 => 8X"70",
        1849 => 8X"1C",
        1850 => 8X"C6",
        1851 => 8X"C6",
        1852 => 8X"7C",
        1853 => 8X"00",
        1854 => 8X"00",
        1855 => 8X"00",
        1856 => 8X"00",
        1857 => 8X"00",
        1858 => 8X"10",
        1859 => 8X"30",
        1860 => 8X"30",
        1861 => 8X"FC",
        1862 => 8X"30",
        1863 => 8X"30",
        1864 => 8X"30",
        1865 => 8X"30",
        1866 => 8X"30",
        1867 => 8X"36",
        1868 => 8X"1C",
        1869 => 8X"00",
        1870 => 8X"00",
        1871 => 8X"00",
        1872 => 8X"00",
        1873 => 8X"00",
        1874 => 8X"00",
        1875 => 8X"00",
        1876 => 8X"00",
        1877 => 8X"CC",
        1878 => 8X"CC",
        1879 => 8X"CC",
        1880 => 8X"CC",
        1881 => 8X"CC",
        1882 => 8X"CC",
        1883 => 8X"CC",
        1884 => 8X"76",
        1885 => 8X"00",
        1886 => 8X"00",
        1887 => 8X"00",
        1888 => 8X"00",
        1889 => 8X"00",
        1890 => 8X"00",
        1891 => 8X"00",
        1892 => 8X"00",
        1893 => 8X"66",
        1894 => 8X"66",
        1895 => 8X"66",
        1896 => 8X"66",
        1897 => 8X"66",
        1898 => 8X"66",
        1899 => 8X"3C",
        1900 => 8X"18",
        1901 => 8X"00",
        1902 => 8X"00",
        1903 => 8X"00",
        1904 => 8X"00",
        1905 => 8X"00",
        1906 => 8X"00",
        1907 => 8X"00",
        1908 => 8X"00",
        1909 => 8X"C6",
        1910 => 8X"C6",
        1911 => 8X"C6",
        1912 => 8X"D6",
        1913 => 8X"D6",
        1914 => 8X"FE",
        1915 => 8X"6C",
        1916 => 8X"6C",
        1917 => 8X"00",
        1918 => 8X"00",
        1919 => 8X"00",
        1920 => 8X"00",
        1921 => 8X"00",
        1922 => 8X"00",
        1923 => 8X"00",
        1924 => 8X"00",
        1925 => 8X"C6",
        1926 => 8X"C6",
        1927 => 8X"6C",
        1928 => 8X"38",
        1929 => 8X"38",
        1930 => 8X"6C",
        1931 => 8X"C6",
        1932 => 8X"C6",
        1933 => 8X"00",
        1934 => 8X"00",
        1935 => 8X"00",
        1936 => 8X"00",
        1937 => 8X"00",
        1938 => 8X"00",
        1939 => 8X"00",
        1940 => 8X"00",
        1941 => 8X"C6",
        1942 => 8X"C6",
        1943 => 8X"C6",
        1944 => 8X"C6",
        1945 => 8X"C6",
        1946 => 8X"C6",
        1947 => 8X"7E",
        1948 => 8X"06",
        1949 => 8X"0C",
        1950 => 8X"F8",
        1951 => 8X"00",
        1952 => 8X"00",
        1953 => 8X"00",
        1954 => 8X"00",
        1955 => 8X"00",
        1956 => 8X"00",
        1957 => 8X"FE",
        1958 => 8X"C6",
        1959 => 8X"CC",
        1960 => 8X"18",
        1961 => 8X"30",
        1962 => 8X"66",
        1963 => 8X"C6",
        1964 => 8X"FE",
        1965 => 8X"00",
        1966 => 8X"00",
        1967 => 8X"00",
        1968 => 8X"00",
        1969 => 8X"0E",
        1970 => 8X"18",
        1971 => 8X"18",
        1972 => 8X"18",
        1973 => 8X"18",
        1974 => 8X"18",
        1975 => 8X"70",
        1976 => 8X"70",
        1977 => 8X"18",
        1978 => 8X"18",
        1979 => 8X"18",
        1980 => 8X"18",
        1981 => 8X"18",
        1982 => 8X"0E",
        1983 => 8X"00",
        1984 => 8X"00",
        1985 => 8X"00",
        1986 => 8X"18",
        1987 => 8X"18",
        1988 => 8X"18",
        1989 => 8X"18",
        1990 => 8X"18",
        1991 => 8X"00",
        1992 => 8X"18",
        1993 => 8X"18",
        1994 => 8X"18",
        1995 => 8X"18",
        1996 => 8X"18",
        1997 => 8X"00",
        1998 => 8X"00",
        1999 => 8X"00",
        2000 => 8X"00",
        2001 => 8X"70",
        2002 => 8X"18",
        2003 => 8X"18",
        2004 => 8X"18",
        2005 => 8X"18",
        2006 => 8X"18",
        2007 => 8X"0E",
        2008 => 8X"0E",
        2009 => 8X"18",
        2010 => 8X"18",
        2011 => 8X"18",
        2012 => 8X"18",
        2013 => 8X"18",
        2014 => 8X"70",
        2015 => 8X"00",
        2016 => 8X"00",
        2017 => 8X"00",
        2018 => 8X"76",
        2019 => 8X"DC",
        2020 => 8X"00",
        2021 => 8X"00",
        2022 => 8X"00",
        2023 => 8X"00",
        2024 => 8X"00",
        2025 => 8X"00",
        2026 => 8X"00",
        2027 => 8X"00",
        2028 => 8X"00",
        2029 => 8X"00",
        2030 => 8X"00",
        2031 => 8X"00",
        2032 => 8X"00",
        2033 => 8X"00",
        2034 => 8X"00",
        2035 => 8X"00",
        2036 => 8X"10",
        2037 => 8X"38",
        2038 => 8X"6C",
        2039 => 8X"C6",
        2040 => 8X"C6",
        2041 => 8X"C6",
        2042 => 8X"C6",
        2043 => 8X"FE",
        2044 => 8X"00",
        2045 => 8X"00",
        2046 => 8X"00",
        2047 => 8X"00",
        2048 => 8X"00",
        2049 => 8X"00",
        2050 => 8X"10",
        2051 => 8X"38",
        2052 => 8X"6C",
        2053 => 8X"C6",
        2054 => 8X"C6",
        2055 => 8X"C6",
        2056 => 8X"FE",
        2057 => 8X"C6",
        2058 => 8X"C6",
        2059 => 8X"C6",
        2060 => 8X"C6",
        2061 => 8X"00",
        2062 => 8X"00",
        2063 => 8X"00",
        2064 => 8X"00",
        2065 => 8X"00",
        2066 => 8X"FE",
        2067 => 8X"66",
        2068 => 8X"62",
        2069 => 8X"60",
        2070 => 8X"7C",
        2071 => 8X"66",
        2072 => 8X"66",
        2073 => 8X"66",
        2074 => 8X"66",
        2075 => 8X"66",
        2076 => 8X"FC",
        2077 => 8X"00",
        2078 => 8X"00",
        2079 => 8X"00",
        2080 => 8X"00",
        2081 => 8X"00",
        2082 => 8X"FC",
        2083 => 8X"66",
        2084 => 8X"66",
        2085 => 8X"66",
        2086 => 8X"7C",
        2087 => 8X"66",
        2088 => 8X"66",
        2089 => 8X"66",
        2090 => 8X"66",
        2091 => 8X"66",
        2092 => 8X"FC",
        2093 => 8X"00",
        2094 => 8X"00",
        2095 => 8X"00",
        2096 => 8X"00",
        2097 => 8X"00",
        2098 => 8X"FE",
        2099 => 8X"66",
        2100 => 8X"62",
        2101 => 8X"60",
        2102 => 8X"60",
        2103 => 8X"60",
        2104 => 8X"60",
        2105 => 8X"60",
        2106 => 8X"60",
        2107 => 8X"60",
        2108 => 8X"F0",
        2109 => 8X"00",
        2110 => 8X"00",
        2111 => 8X"00",
        2112 => 8X"00",
        2113 => 8X"00",
        2114 => 8X"3E",
        2115 => 8X"66",
        2116 => 8X"66",
        2117 => 8X"66",
        2118 => 8X"66",
        2119 => 8X"66",
        2120 => 8X"66",
        2121 => 8X"66",
        2122 => 8X"66",
        2123 => 8X"66",
        2124 => 8X"FF",
        2125 => 8X"C3",
        2126 => 8X"C3",
        2127 => 8X"00",
        2128 => 8X"00",
        2129 => 8X"00",
        2130 => 8X"FE",
        2131 => 8X"66",
        2132 => 8X"66",
        2133 => 8X"62",
        2134 => 8X"68",
        2135 => 8X"78",
        2136 => 8X"68",
        2137 => 8X"62",
        2138 => 8X"66",
        2139 => 8X"66",
        2140 => 8X"FE",
        2141 => 8X"00",
        2142 => 8X"00",
        2143 => 8X"00",
        2144 => 8X"00",
        2145 => 8X"00",
        2146 => 8X"D6",
        2147 => 8X"D6",
        2148 => 8X"D6",
        2149 => 8X"7C",
        2150 => 8X"38",
        2151 => 8X"7C",
        2152 => 8X"D6",
        2153 => 8X"D6",
        2154 => 8X"D6",
        2155 => 8X"D6",
        2156 => 8X"D6",
        2157 => 8X"00",
        2158 => 8X"00",
        2159 => 8X"00",
        2160 => 8X"00",
        2161 => 8X"00",
        2162 => 8X"7C",
        2163 => 8X"C6",
        2164 => 8X"06",
        2165 => 8X"06",
        2166 => 8X"06",
        2167 => 8X"3C",
        2168 => 8X"06",
        2169 => 8X"06",
        2170 => 8X"06",
        2171 => 8X"C6",
        2172 => 8X"7C",
        2173 => 8X"00",
        2174 => 8X"00",
        2175 => 8X"00",
        2176 => 8X"00",
        2177 => 8X"00",
        2178 => 8X"C6",
        2179 => 8X"C6",
        2180 => 8X"CE",
        2181 => 8X"DE",
        2182 => 8X"FE",
        2183 => 8X"F6",
        2184 => 8X"E6",
        2185 => 8X"C6",
        2186 => 8X"C6",
        2187 => 8X"C6",
        2188 => 8X"C6",
        2189 => 8X"00",
        2190 => 8X"00",
        2191 => 8X"00",
        2192 => 8X"38",
        2193 => 8X"38",
        2194 => 8X"C6",
        2195 => 8X"C6",
        2196 => 8X"CE",
        2197 => 8X"DE",
        2198 => 8X"FE",
        2199 => 8X"F6",
        2200 => 8X"E6",
        2201 => 8X"C6",
        2202 => 8X"C6",
        2203 => 8X"C6",
        2204 => 8X"C6",
        2205 => 8X"00",
        2206 => 8X"00",
        2207 => 8X"00",
        2208 => 8X"00",
        2209 => 8X"00",
        2210 => 8X"E6",
        2211 => 8X"66",
        2212 => 8X"6C",
        2213 => 8X"6C",
        2214 => 8X"78",
        2215 => 8X"6C",
        2216 => 8X"6C",
        2217 => 8X"66",
        2218 => 8X"66",
        2219 => 8X"66",
        2220 => 8X"E6",
        2221 => 8X"00",
        2222 => 8X"00",
        2223 => 8X"00",
        2224 => 8X"00",
        2225 => 8X"00",
        2226 => 8X"3E",
        2227 => 8X"66",
        2228 => 8X"66",
        2229 => 8X"66",
        2230 => 8X"66",
        2231 => 8X"66",
        2232 => 8X"66",
        2233 => 8X"66",
        2234 => 8X"66",
        2235 => 8X"66",
        2236 => 8X"E6",
        2237 => 8X"00",
        2238 => 8X"00",
        2239 => 8X"00",
        2240 => 8X"00",
        2241 => 8X"00",
        2242 => 8X"C6",
        2243 => 8X"EE",
        2244 => 8X"FE",
        2245 => 8X"FE",
        2246 => 8X"D6",
        2247 => 8X"C6",
        2248 => 8X"C6",
        2249 => 8X"C6",
        2250 => 8X"C6",
        2251 => 8X"C6",
        2252 => 8X"C6",
        2253 => 8X"00",
        2254 => 8X"00",
        2255 => 8X"00",
        2256 => 8X"00",
        2257 => 8X"00",
        2258 => 8X"C6",
        2259 => 8X"C6",
        2260 => 8X"C6",
        2261 => 8X"C6",
        2262 => 8X"FE",
        2263 => 8X"C6",
        2264 => 8X"C6",
        2265 => 8X"C6",
        2266 => 8X"C6",
        2267 => 8X"C6",
        2268 => 8X"C6",
        2269 => 8X"00",
        2270 => 8X"00",
        2271 => 8X"00",
        2272 => 8X"00",
        2273 => 8X"00",
        2274 => 8X"7C",
        2275 => 8X"C6",
        2276 => 8X"C6",
        2277 => 8X"C6",
        2278 => 8X"C6",
        2279 => 8X"C6",
        2280 => 8X"C6",
        2281 => 8X"C6",
        2282 => 8X"C6",
        2283 => 8X"C6",
        2284 => 8X"7C",
        2285 => 8X"00",
        2286 => 8X"00",
        2287 => 8X"00",
        2288 => 8X"00",
        2289 => 8X"00",
        2290 => 8X"FE",
        2291 => 8X"C6",
        2292 => 8X"C6",
        2293 => 8X"C6",
        2294 => 8X"C6",
        2295 => 8X"C6",
        2296 => 8X"C6",
        2297 => 8X"C6",
        2298 => 8X"C6",
        2299 => 8X"C6",
        2300 => 8X"C6",
        2301 => 8X"00",
        2302 => 8X"00",
        2303 => 8X"00",
        2304 => 8X"00",
        2305 => 8X"00",
        2306 => 8X"FC",
        2307 => 8X"66",
        2308 => 8X"66",
        2309 => 8X"66",
        2310 => 8X"66",
        2311 => 8X"66",
        2312 => 8X"7C",
        2313 => 8X"60",
        2314 => 8X"60",
        2315 => 8X"60",
        2316 => 8X"F0",
        2317 => 8X"00",
        2318 => 8X"00",
        2319 => 8X"00",
        2320 => 8X"00",
        2321 => 8X"00",
        2322 => 8X"7C",
        2323 => 8X"C6",
        2324 => 8X"C6",
        2325 => 8X"C0",
        2326 => 8X"C0",
        2327 => 8X"C0",
        2328 => 8X"C0",
        2329 => 8X"C6",
        2330 => 8X"C6",
        2331 => 8X"C6",
        2332 => 8X"7C",
        2333 => 8X"00",
        2334 => 8X"00",
        2335 => 8X"00",
        2336 => 8X"00",
        2337 => 8X"00",
        2338 => 8X"7E",
        2339 => 8X"7E",
        2340 => 8X"5A",
        2341 => 8X"18",
        2342 => 8X"18",
        2343 => 8X"18",
        2344 => 8X"18",
        2345 => 8X"18",
        2346 => 8X"18",
        2347 => 8X"18",
        2348 => 8X"3C",
        2349 => 8X"00",
        2350 => 8X"00",
        2351 => 8X"00",
        2352 => 8X"00",
        2353 => 8X"00",
        2354 => 8X"C6",
        2355 => 8X"C6",
        2356 => 8X"C6",
        2357 => 8X"C6",
        2358 => 8X"C6",
        2359 => 8X"7E",
        2360 => 8X"06",
        2361 => 8X"06",
        2362 => 8X"06",
        2363 => 8X"C6",
        2364 => 8X"7C",
        2365 => 8X"00",
        2366 => 8X"00",
        2367 => 8X"00",
        2368 => 8X"00",
        2369 => 8X"00",
        2370 => 8X"18",
        2371 => 8X"7E",
        2372 => 8X"DB",
        2373 => 8X"DB",
        2374 => 8X"DB",
        2375 => 8X"DB",
        2376 => 8X"DB",
        2377 => 8X"DB",
        2378 => 8X"DB",
        2379 => 8X"7E",
        2380 => 8X"18",
        2381 => 8X"00",
        2382 => 8X"00",
        2383 => 8X"00",
        2384 => 8X"00",
        2385 => 8X"00",
        2386 => 8X"C6",
        2387 => 8X"C6",
        2388 => 8X"C6",
        2389 => 8X"6C",
        2390 => 8X"38",
        2391 => 8X"38",
        2392 => 8X"38",
        2393 => 8X"6C",
        2394 => 8X"C6",
        2395 => 8X"C6",
        2396 => 8X"C6",
        2397 => 8X"00",
        2398 => 8X"00",
        2399 => 8X"00",
        2400 => 8X"00",
        2401 => 8X"00",
        2402 => 8X"CC",
        2403 => 8X"CC",
        2404 => 8X"CC",
        2405 => 8X"CC",
        2406 => 8X"CC",
        2407 => 8X"CC",
        2408 => 8X"CC",
        2409 => 8X"CC",
        2410 => 8X"CC",
        2411 => 8X"CC",
        2412 => 8X"FE",
        2413 => 8X"06",
        2414 => 8X"06",
        2415 => 8X"00",
        2416 => 8X"00",
        2417 => 8X"00",
        2418 => 8X"C6",
        2419 => 8X"C6",
        2420 => 8X"C6",
        2421 => 8X"C6",
        2422 => 8X"C6",
        2423 => 8X"C6",
        2424 => 8X"7E",
        2425 => 8X"06",
        2426 => 8X"06",
        2427 => 8X"06",
        2428 => 8X"06",
        2429 => 8X"00",
        2430 => 8X"00",
        2431 => 8X"00",
        2432 => 8X"00",
        2433 => 8X"00",
        2434 => 8X"D6",
        2435 => 8X"D6",
        2436 => 8X"D6",
        2437 => 8X"D6",
        2438 => 8X"D6",
        2439 => 8X"D6",
        2440 => 8X"D6",
        2441 => 8X"D6",
        2442 => 8X"D6",
        2443 => 8X"D6",
        2444 => 8X"FE",
        2445 => 8X"00",
        2446 => 8X"00",
        2447 => 8X"00",
        2448 => 8X"00",
        2449 => 8X"00",
        2450 => 8X"D6",
        2451 => 8X"D6",
        2452 => 8X"D6",
        2453 => 8X"D6",
        2454 => 8X"D6",
        2455 => 8X"D6",
        2456 => 8X"D6",
        2457 => 8X"D6",
        2458 => 8X"D6",
        2459 => 8X"D6",
        2460 => 8X"FE",
        2461 => 8X"03",
        2462 => 8X"03",
        2463 => 8X"00",
        2464 => 8X"00",
        2465 => 8X"00",
        2466 => 8X"F8",
        2467 => 8X"F0",
        2468 => 8X"B0",
        2469 => 8X"30",
        2470 => 8X"3C",
        2471 => 8X"36",
        2472 => 8X"36",
        2473 => 8X"36",
        2474 => 8X"36",
        2475 => 8X"36",
        2476 => 8X"7C",
        2477 => 8X"00",
        2478 => 8X"00",
        2479 => 8X"00",
        2480 => 8X"00",
        2481 => 8X"00",
        2482 => 8X"C6",
        2483 => 8X"C6",
        2484 => 8X"C6",
        2485 => 8X"C6",
        2486 => 8X"F6",
        2487 => 8X"DE",
        2488 => 8X"DE",
        2489 => 8X"DE",
        2490 => 8X"DE",
        2491 => 8X"DE",
        2492 => 8X"F6",
        2493 => 8X"00",
        2494 => 8X"00",
        2495 => 8X"00",
        2496 => 8X"00",
        2497 => 8X"00",
        2498 => 8X"F0",
        2499 => 8X"60",
        2500 => 8X"60",
        2501 => 8X"60",
        2502 => 8X"7C",
        2503 => 8X"66",
        2504 => 8X"66",
        2505 => 8X"66",
        2506 => 8X"66",
        2507 => 8X"66",
        2508 => 8X"FC",
        2509 => 8X"00",
        2510 => 8X"00",
        2511 => 8X"00",
        2512 => 8X"00",
        2513 => 8X"00",
        2514 => 8X"78",
        2515 => 8X"CC",
        2516 => 8X"86",
        2517 => 8X"86",
        2518 => 8X"26",
        2519 => 8X"3E",
        2520 => 8X"26",
        2521 => 8X"86",
        2522 => 8X"86",
        2523 => 8X"CC",
        2524 => 8X"78",
        2525 => 8X"00",
        2526 => 8X"00",
        2527 => 8X"00",
        2528 => 8X"00",
        2529 => 8X"00",
        2530 => 8X"9C",
        2531 => 8X"B6",
        2532 => 8X"B6",
        2533 => 8X"B6",
        2534 => 8X"B6",
        2535 => 8X"F6",
        2536 => 8X"B6",
        2537 => 8X"B6",
        2538 => 8X"B6",
        2539 => 8X"B6",
        2540 => 8X"9C",
        2541 => 8X"00",
        2542 => 8X"00",
        2543 => 8X"00",
        2544 => 8X"00",
        2545 => 8X"00",
        2546 => 8X"7E",
        2547 => 8X"CC",
        2548 => 8X"CC",
        2549 => 8X"CC",
        2550 => 8X"CC",
        2551 => 8X"7C",
        2552 => 8X"6C",
        2553 => 8X"CC",
        2554 => 8X"CC",
        2555 => 8X"CE",
        2556 => 8X"CE",
        2557 => 8X"00",
        2558 => 8X"00",
        2559 => 8X"00",
        2560 => 8X"00",
        2561 => 8X"00",
        2562 => 8X"00",
        2563 => 8X"00",
        2564 => 8X"00",
        2565 => 8X"78",
        2566 => 8X"CC",
        2567 => 8X"0C",
        2568 => 8X"7C",
        2569 => 8X"CC",
        2570 => 8X"CC",
        2571 => 8X"CC",
        2572 => 8X"76",
        2573 => 8X"00",
        2574 => 8X"00",
        2575 => 8X"00",
        2576 => 8X"00",
        2577 => 8X"00",
        2578 => 8X"00",
        2579 => 8X"1C",
        2580 => 8X"30",
        2581 => 8X"60",
        2582 => 8X"7C",
        2583 => 8X"66",
        2584 => 8X"66",
        2585 => 8X"66",
        2586 => 8X"66",
        2587 => 8X"66",
        2588 => 8X"3C",
        2589 => 8X"00",
        2590 => 8X"00",
        2591 => 8X"00",
        2592 => 8X"00",
        2593 => 8X"00",
        2594 => 8X"00",
        2595 => 8X"00",
        2596 => 8X"00",
        2597 => 8X"FC",
        2598 => 8X"66",
        2599 => 8X"66",
        2600 => 8X"7C",
        2601 => 8X"66",
        2602 => 8X"66",
        2603 => 8X"66",
        2604 => 8X"FC",
        2605 => 8X"00",
        2606 => 8X"00",
        2607 => 8X"00",
        2608 => 8X"00",
        2609 => 8X"00",
        2610 => 8X"00",
        2611 => 8X"00",
        2612 => 8X"00",
        2613 => 8X"FE",
        2614 => 8X"62",
        2615 => 8X"60",
        2616 => 8X"60",
        2617 => 8X"60",
        2618 => 8X"60",
        2619 => 8X"60",
        2620 => 8X"F0",
        2621 => 8X"00",
        2622 => 8X"00",
        2623 => 8X"00",
        2624 => 8X"00",
        2625 => 8X"00",
        2626 => 8X"00",
        2627 => 8X"00",
        2628 => 8X"00",
        2629 => 8X"3E",
        2630 => 8X"66",
        2631 => 8X"66",
        2632 => 8X"66",
        2633 => 8X"66",
        2634 => 8X"66",
        2635 => 8X"66",
        2636 => 8X"FF",
        2637 => 8X"C3",
        2638 => 8X"C3",
        2639 => 8X"00",
        2640 => 8X"00",
        2641 => 8X"00",
        2642 => 8X"00",
        2643 => 8X"00",
        2644 => 8X"00",
        2645 => 8X"7C",
        2646 => 8X"C6",
        2647 => 8X"C6",
        2648 => 8X"FE",
        2649 => 8X"C0",
        2650 => 8X"C0",
        2651 => 8X"C6",
        2652 => 8X"7C",
        2653 => 8X"00",
        2654 => 8X"00",
        2655 => 8X"00",
        2656 => 8X"00",
        2657 => 8X"00",
        2658 => 8X"00",
        2659 => 8X"00",
        2660 => 8X"00",
        2661 => 8X"D6",
        2662 => 8X"D6",
        2663 => 8X"D6",
        2664 => 8X"7C",
        2665 => 8X"7C",
        2666 => 8X"D6",
        2667 => 8X"D6",
        2668 => 8X"D6",
        2669 => 8X"00",
        2670 => 8X"00",
        2671 => 8X"00",
        2672 => 8X"00",
        2673 => 8X"00",
        2674 => 8X"00",
        2675 => 8X"00",
        2676 => 8X"00",
        2677 => 8X"3C",
        2678 => 8X"66",
        2679 => 8X"66",
        2680 => 8X"0C",
        2681 => 8X"06",
        2682 => 8X"66",
        2683 => 8X"66",
        2684 => 8X"3C",
        2685 => 8X"00",
        2686 => 8X"00",
        2687 => 8X"00",
        2688 => 8X"00",
        2689 => 8X"00",
        2690 => 8X"00",
        2691 => 8X"00",
        2692 => 8X"00",
        2693 => 8X"C6",
        2694 => 8X"CE",
        2695 => 8X"DE",
        2696 => 8X"FE",
        2697 => 8X"F6",
        2698 => 8X"E6",
        2699 => 8X"C6",
        2700 => 8X"C6",
        2701 => 8X"00",
        2702 => 8X"00",
        2703 => 8X"00",
        2704 => 8X"00",
        2705 => 8X"00",
        2706 => 8X"38",
        2707 => 8X"38",
        2708 => 8X"00",
        2709 => 8X"C6",
        2710 => 8X"CE",
        2711 => 8X"DE",
        2712 => 8X"FE",
        2713 => 8X"F6",
        2714 => 8X"E6",
        2715 => 8X"C6",
        2716 => 8X"C6",
        2717 => 8X"00",
        2718 => 8X"00",
        2719 => 8X"00",
        2720 => 8X"00",
        2721 => 8X"00",
        2722 => 8X"00",
        2723 => 8X"00",
        2724 => 8X"00",
        2725 => 8X"E6",
        2726 => 8X"66",
        2727 => 8X"6C",
        2728 => 8X"78",
        2729 => 8X"6C",
        2730 => 8X"66",
        2731 => 8X"66",
        2732 => 8X"E6",
        2733 => 8X"00",
        2734 => 8X"00",
        2735 => 8X"00",
        2736 => 8X"00",
        2737 => 8X"00",
        2738 => 8X"00",
        2739 => 8X"00",
        2740 => 8X"00",
        2741 => 8X"3E",
        2742 => 8X"66",
        2743 => 8X"66",
        2744 => 8X"66",
        2745 => 8X"66",
        2746 => 8X"66",
        2747 => 8X"66",
        2748 => 8X"E6",
        2749 => 8X"00",
        2750 => 8X"00",
        2751 => 8X"00",
        2752 => 8X"00",
        2753 => 8X"00",
        2754 => 8X"00",
        2755 => 8X"00",
        2756 => 8X"00",
        2757 => 8X"C6",
        2758 => 8X"EE",
        2759 => 8X"FE",
        2760 => 8X"FE",
        2761 => 8X"D6",
        2762 => 8X"C6",
        2763 => 8X"C6",
        2764 => 8X"C6",
        2765 => 8X"00",
        2766 => 8X"00",
        2767 => 8X"00",
        2768 => 8X"00",
        2769 => 8X"00",
        2770 => 8X"00",
        2771 => 8X"00",
        2772 => 8X"00",
        2773 => 8X"C6",
        2774 => 8X"C6",
        2775 => 8X"C6",
        2776 => 8X"FE",
        2777 => 8X"C6",
        2778 => 8X"C6",
        2779 => 8X"C6",
        2780 => 8X"C6",
        2781 => 8X"00",
        2782 => 8X"00",
        2783 => 8X"00",
        2784 => 8X"00",
        2785 => 8X"00",
        2786 => 8X"00",
        2787 => 8X"00",
        2788 => 8X"00",
        2789 => 8X"7C",
        2790 => 8X"C6",
        2791 => 8X"C6",
        2792 => 8X"C6",
        2793 => 8X"C6",
        2794 => 8X"C6",
        2795 => 8X"C6",
        2796 => 8X"7C",
        2797 => 8X"00",
        2798 => 8X"00",
        2799 => 8X"00",
        2800 => 8X"00",
        2801 => 8X"00",
        2802 => 8X"00",
        2803 => 8X"00",
        2804 => 8X"00",
        2805 => 8X"FE",
        2806 => 8X"C6",
        2807 => 8X"C6",
        2808 => 8X"C6",
        2809 => 8X"C6",
        2810 => 8X"C6",
        2811 => 8X"C6",
        2812 => 8X"C6",
        2813 => 8X"00",
        2814 => 8X"00",
        2815 => 8X"00",
        2816 => 8X"44",
        2817 => 8X"11",
        2818 => 8X"44",
        2819 => 8X"11",
        2820 => 8X"44",
        2821 => 8X"11",
        2822 => 8X"44",
        2823 => 8X"11",
        2824 => 8X"44",
        2825 => 8X"11",
        2826 => 8X"44",
        2827 => 8X"11",
        2828 => 8X"44",
        2829 => 8X"11",
        2830 => 8X"44",
        2831 => 8X"11",
        2832 => 8X"AA",
        2833 => 8X"55",
        2834 => 8X"AA",
        2835 => 8X"55",
        2836 => 8X"AA",
        2837 => 8X"55",
        2838 => 8X"AA",
        2839 => 8X"55",
        2840 => 8X"AA",
        2841 => 8X"55",
        2842 => 8X"AA",
        2843 => 8X"55",
        2844 => 8X"AA",
        2845 => 8X"55",
        2846 => 8X"AA",
        2847 => 8X"55",
        2848 => 8X"77",
        2849 => 8X"DD",
        2850 => 8X"77",
        2851 => 8X"DD",
        2852 => 8X"77",
        2853 => 8X"DD",
        2854 => 8X"77",
        2855 => 8X"DD",
        2856 => 8X"77",
        2857 => 8X"DD",
        2858 => 8X"77",
        2859 => 8X"DD",
        2860 => 8X"77",
        2861 => 8X"DD",
        2862 => 8X"77",
        2863 => 8X"DD",
        2864 => 8X"18",
        2865 => 8X"18",
        2866 => 8X"18",
        2867 => 8X"18",
        2868 => 8X"18",
        2869 => 8X"18",
        2870 => 8X"18",
        2871 => 8X"18",
        2872 => 8X"18",
        2873 => 8X"18",
        2874 => 8X"18",
        2875 => 8X"18",
        2876 => 8X"18",
        2877 => 8X"18",
        2878 => 8X"18",
        2879 => 8X"18",
        2880 => 8X"18",
        2881 => 8X"18",
        2882 => 8X"18",
        2883 => 8X"18",
        2884 => 8X"18",
        2885 => 8X"18",
        2886 => 8X"18",
        2887 => 8X"18",
        2888 => 8X"F8",
        2889 => 8X"18",
        2890 => 8X"18",
        2891 => 8X"18",
        2892 => 8X"18",
        2893 => 8X"18",
        2894 => 8X"18",
        2895 => 8X"18",
        2896 => 8X"18",
        2897 => 8X"18",
        2898 => 8X"18",
        2899 => 8X"18",
        2900 => 8X"18",
        2901 => 8X"18",
        2902 => 8X"F8",
        2903 => 8X"18",
        2904 => 8X"F8",
        2905 => 8X"18",
        2906 => 8X"18",
        2907 => 8X"18",
        2908 => 8X"18",
        2909 => 8X"18",
        2910 => 8X"18",
        2911 => 8X"18",
        2912 => 8X"36",
        2913 => 8X"36",
        2914 => 8X"36",
        2915 => 8X"36",
        2916 => 8X"36",
        2917 => 8X"36",
        2918 => 8X"36",
        2919 => 8X"36",
        2920 => 8X"F6",
        2921 => 8X"36",
        2922 => 8X"36",
        2923 => 8X"36",
        2924 => 8X"36",
        2925 => 8X"36",
        2926 => 8X"36",
        2927 => 8X"36",
        2928 => 8X"00",
        2929 => 8X"00",
        2930 => 8X"00",
        2931 => 8X"00",
        2932 => 8X"00",
        2933 => 8X"00",
        2934 => 8X"00",
        2935 => 8X"00",
        2936 => 8X"FE",
        2937 => 8X"36",
        2938 => 8X"36",
        2939 => 8X"36",
        2940 => 8X"36",
        2941 => 8X"36",
        2942 => 8X"36",
        2943 => 8X"36",
        2944 => 8X"00",
        2945 => 8X"00",
        2946 => 8X"00",
        2947 => 8X"00",
        2948 => 8X"00",
        2949 => 8X"00",
        2950 => 8X"F8",
        2951 => 8X"18",
        2952 => 8X"F8",
        2953 => 8X"18",
        2954 => 8X"18",
        2955 => 8X"18",
        2956 => 8X"18",
        2957 => 8X"18",
        2958 => 8X"18",
        2959 => 8X"18",
        2960 => 8X"36",
        2961 => 8X"36",
        2962 => 8X"36",
        2963 => 8X"36",
        2964 => 8X"36",
        2965 => 8X"36",
        2966 => 8X"F6",
        2967 => 8X"06",
        2968 => 8X"F6",
        2969 => 8X"36",
        2970 => 8X"36",
        2971 => 8X"36",
        2972 => 8X"36",
        2973 => 8X"36",
        2974 => 8X"36",
        2975 => 8X"36",
        2976 => 8X"36",
        2977 => 8X"36",
        2978 => 8X"36",
        2979 => 8X"36",
        2980 => 8X"36",
        2981 => 8X"36",
        2982 => 8X"36",
        2983 => 8X"36",
        2984 => 8X"36",
        2985 => 8X"36",
        2986 => 8X"36",
        2987 => 8X"36",
        2988 => 8X"36",
        2989 => 8X"36",
        2990 => 8X"36",
        2991 => 8X"36",
        2992 => 8X"00",
        2993 => 8X"00",
        2994 => 8X"00",
        2995 => 8X"00",
        2996 => 8X"00",
        2997 => 8X"00",
        2998 => 8X"FE",
        2999 => 8X"06",
        3000 => 8X"F6",
        3001 => 8X"36",
        3002 => 8X"36",
        3003 => 8X"36",
        3004 => 8X"36",
        3005 => 8X"36",
        3006 => 8X"36",
        3007 => 8X"36",
        3008 => 8X"36",
        3009 => 8X"36",
        3010 => 8X"36",
        3011 => 8X"36",
        3012 => 8X"36",
        3013 => 8X"36",
        3014 => 8X"F6",
        3015 => 8X"06",
        3016 => 8X"FE",
        3017 => 8X"00",
        3018 => 8X"00",
        3019 => 8X"00",
        3020 => 8X"00",
        3021 => 8X"00",
        3022 => 8X"00",
        3023 => 8X"00",
        3024 => 8X"36",
        3025 => 8X"36",
        3026 => 8X"36",
        3027 => 8X"36",
        3028 => 8X"36",
        3029 => 8X"36",
        3030 => 8X"36",
        3031 => 8X"36",
        3032 => 8X"FE",
        3033 => 8X"00",
        3034 => 8X"00",
        3035 => 8X"00",
        3036 => 8X"00",
        3037 => 8X"00",
        3038 => 8X"00",
        3039 => 8X"00",
        3040 => 8X"18",
        3041 => 8X"18",
        3042 => 8X"18",
        3043 => 8X"18",
        3044 => 8X"18",
        3045 => 8X"18",
        3046 => 8X"F8",
        3047 => 8X"18",
        3048 => 8X"F8",
        3049 => 8X"00",
        3050 => 8X"00",
        3051 => 8X"00",
        3052 => 8X"00",
        3053 => 8X"00",
        3054 => 8X"00",
        3055 => 8X"00",
        3056 => 8X"00",
        3057 => 8X"00",
        3058 => 8X"00",
        3059 => 8X"00",
        3060 => 8X"00",
        3061 => 8X"00",
        3062 => 8X"00",
        3063 => 8X"00",
        3064 => 8X"F8",
        3065 => 8X"18",
        3066 => 8X"18",
        3067 => 8X"18",
        3068 => 8X"18",
        3069 => 8X"18",
        3070 => 8X"18",
        3071 => 8X"18",
        3072 => 8X"18",
        3073 => 8X"18",
        3074 => 8X"18",
        3075 => 8X"18",
        3076 => 8X"18",
        3077 => 8X"18",
        3078 => 8X"18",
        3079 => 8X"18",
        3080 => 8X"1F",
        3081 => 8X"00",
        3082 => 8X"00",
        3083 => 8X"00",
        3084 => 8X"00",
        3085 => 8X"00",
        3086 => 8X"00",
        3087 => 8X"00",
        3088 => 8X"18",
        3089 => 8X"18",
        3090 => 8X"18",
        3091 => 8X"18",
        3092 => 8X"18",
        3093 => 8X"18",
        3094 => 8X"18",
        3095 => 8X"18",
        3096 => 8X"FF",
        3097 => 8X"00",
        3098 => 8X"00",
        3099 => 8X"00",
        3100 => 8X"00",
        3101 => 8X"00",
        3102 => 8X"00",
        3103 => 8X"00",
        3104 => 8X"00",
        3105 => 8X"00",
        3106 => 8X"00",
        3107 => 8X"00",
        3108 => 8X"00",
        3109 => 8X"00",
        3110 => 8X"00",
        3111 => 8X"00",
        3112 => 8X"FF",
        3113 => 8X"18",
        3114 => 8X"18",
        3115 => 8X"18",
        3116 => 8X"18",
        3117 => 8X"18",
        3118 => 8X"18",
        3119 => 8X"18",
        3120 => 8X"18",
        3121 => 8X"18",
        3122 => 8X"18",
        3123 => 8X"18",
        3124 => 8X"18",
        3125 => 8X"18",
        3126 => 8X"18",
        3127 => 8X"18",
        3128 => 8X"1F",
        3129 => 8X"18",
        3130 => 8X"18",
        3131 => 8X"18",
        3132 => 8X"18",
        3133 => 8X"18",
        3134 => 8X"18",
        3135 => 8X"18",
        3136 => 8X"00",
        3137 => 8X"00",
        3138 => 8X"00",
        3139 => 8X"00",
        3140 => 8X"00",
        3141 => 8X"00",
        3142 => 8X"00",
        3143 => 8X"00",
        3144 => 8X"FF",
        3145 => 8X"00",
        3146 => 8X"00",
        3147 => 8X"00",
        3148 => 8X"00",
        3149 => 8X"00",
        3150 => 8X"00",
        3151 => 8X"00",
        3152 => 8X"18",
        3153 => 8X"18",
        3154 => 8X"18",
        3155 => 8X"18",
        3156 => 8X"18",
        3157 => 8X"18",
        3158 => 8X"18",
        3159 => 8X"18",
        3160 => 8X"FF",
        3161 => 8X"18",
        3162 => 8X"18",
        3163 => 8X"18",
        3164 => 8X"18",
        3165 => 8X"18",
        3166 => 8X"18",
        3167 => 8X"18",
        3168 => 8X"18",
        3169 => 8X"18",
        3170 => 8X"18",
        3171 => 8X"18",
        3172 => 8X"18",
        3173 => 8X"18",
        3174 => 8X"1F",
        3175 => 8X"18",
        3176 => 8X"1F",
        3177 => 8X"18",
        3178 => 8X"18",
        3179 => 8X"18",
        3180 => 8X"18",
        3181 => 8X"18",
        3182 => 8X"18",
        3183 => 8X"18",
        3184 => 8X"36",
        3185 => 8X"36",
        3186 => 8X"36",
        3187 => 8X"36",
        3188 => 8X"36",
        3189 => 8X"36",
        3190 => 8X"36",
        3191 => 8X"36",
        3192 => 8X"37",
        3193 => 8X"36",
        3194 => 8X"36",
        3195 => 8X"36",
        3196 => 8X"36",
        3197 => 8X"36",
        3198 => 8X"36",
        3199 => 8X"36",
        3200 => 8X"36",
        3201 => 8X"36",
        3202 => 8X"36",
        3203 => 8X"36",
        3204 => 8X"36",
        3205 => 8X"36",
        3206 => 8X"37",
        3207 => 8X"30",
        3208 => 8X"3F",
        3209 => 8X"00",
        3210 => 8X"00",
        3211 => 8X"00",
        3212 => 8X"00",
        3213 => 8X"00",
        3214 => 8X"00",
        3215 => 8X"00",
        3216 => 8X"00",
        3217 => 8X"00",
        3218 => 8X"00",
        3219 => 8X"00",
        3220 => 8X"00",
        3221 => 8X"00",
        3222 => 8X"3F",
        3223 => 8X"30",
        3224 => 8X"37",
        3225 => 8X"36",
        3226 => 8X"36",
        3227 => 8X"36",
        3228 => 8X"36",
        3229 => 8X"36",
        3230 => 8X"36",
        3231 => 8X"36",
        3232 => 8X"36",
        3233 => 8X"36",
        3234 => 8X"36",
        3235 => 8X"36",
        3236 => 8X"36",
        3237 => 8X"36",
        3238 => 8X"F7",
        3239 => 8X"00",
        3240 => 8X"FF",
        3241 => 8X"00",
        3242 => 8X"00",
        3243 => 8X"00",
        3244 => 8X"00",
        3245 => 8X"00",
        3246 => 8X"00",
        3247 => 8X"00",
        3248 => 8X"00",
        3249 => 8X"00",
        3250 => 8X"00",
        3251 => 8X"00",
        3252 => 8X"00",
        3253 => 8X"00",
        3254 => 8X"FF",
        3255 => 8X"00",
        3256 => 8X"F7",
        3257 => 8X"36",
        3258 => 8X"36",
        3259 => 8X"36",
        3260 => 8X"36",
        3261 => 8X"36",
        3262 => 8X"36",
        3263 => 8X"36",
        3264 => 8X"36",
        3265 => 8X"36",
        3266 => 8X"36",
        3267 => 8X"36",
        3268 => 8X"36",
        3269 => 8X"36",
        3270 => 8X"37",
        3271 => 8X"30",
        3272 => 8X"37",
        3273 => 8X"36",
        3274 => 8X"36",
        3275 => 8X"36",
        3276 => 8X"36",
        3277 => 8X"36",
        3278 => 8X"36",
        3279 => 8X"36",
        3280 => 8X"00",
        3281 => 8X"00",
        3282 => 8X"00",
        3283 => 8X"00",
        3284 => 8X"00",
        3285 => 8X"00",
        3286 => 8X"FF",
        3287 => 8X"00",
        3288 => 8X"FF",
        3289 => 8X"00",
        3290 => 8X"00",
        3291 => 8X"00",
        3292 => 8X"00",
        3293 => 8X"00",
        3294 => 8X"00",
        3295 => 8X"00",
        3296 => 8X"36",
        3297 => 8X"36",
        3298 => 8X"36",
        3299 => 8X"36",
        3300 => 8X"36",
        3301 => 8X"36",
        3302 => 8X"F7",
        3303 => 8X"00",
        3304 => 8X"F7",
        3305 => 8X"36",
        3306 => 8X"36",
        3307 => 8X"36",
        3308 => 8X"36",
        3309 => 8X"36",
        3310 => 8X"36",
        3311 => 8X"36",
        3312 => 8X"18",
        3313 => 8X"18",
        3314 => 8X"18",
        3315 => 8X"18",
        3316 => 8X"18",
        3317 => 8X"18",
        3318 => 8X"FF",
        3319 => 8X"00",
        3320 => 8X"FF",
        3321 => 8X"00",
        3322 => 8X"00",
        3323 => 8X"00",
        3324 => 8X"00",
        3325 => 8X"00",
        3326 => 8X"00",
        3327 => 8X"00",
        3328 => 8X"36",
        3329 => 8X"36",
        3330 => 8X"36",
        3331 => 8X"36",
        3332 => 8X"36",
        3333 => 8X"36",
        3334 => 8X"36",
        3335 => 8X"36",
        3336 => 8X"FF",
        3337 => 8X"00",
        3338 => 8X"00",
        3339 => 8X"00",
        3340 => 8X"00",
        3341 => 8X"00",
        3342 => 8X"00",
        3343 => 8X"00",
        3344 => 8X"00",
        3345 => 8X"00",
        3346 => 8X"00",
        3347 => 8X"00",
        3348 => 8X"00",
        3349 => 8X"00",
        3350 => 8X"FF",
        3351 => 8X"00",
        3352 => 8X"FF",
        3353 => 8X"18",
        3354 => 8X"18",
        3355 => 8X"18",
        3356 => 8X"18",
        3357 => 8X"18",
        3358 => 8X"18",
        3359 => 8X"18",
        3360 => 8X"00",
        3361 => 8X"00",
        3362 => 8X"00",
        3363 => 8X"00",
        3364 => 8X"00",
        3365 => 8X"00",
        3366 => 8X"00",
        3367 => 8X"00",
        3368 => 8X"FF",
        3369 => 8X"36",
        3370 => 8X"36",
        3371 => 8X"36",
        3372 => 8X"36",
        3373 => 8X"36",
        3374 => 8X"36",
        3375 => 8X"36",
        3376 => 8X"36",
        3377 => 8X"36",
        3378 => 8X"36",
        3379 => 8X"36",
        3380 => 8X"36",
        3381 => 8X"36",
        3382 => 8X"36",
        3383 => 8X"36",
        3384 => 8X"3F",
        3385 => 8X"00",
        3386 => 8X"00",
        3387 => 8X"00",
        3388 => 8X"00",
        3389 => 8X"00",
        3390 => 8X"00",
        3391 => 8X"00",
        3392 => 8X"18",
        3393 => 8X"18",
        3394 => 8X"18",
        3395 => 8X"18",
        3396 => 8X"18",
        3397 => 8X"18",
        3398 => 8X"1F",
        3399 => 8X"18",
        3400 => 8X"1F",
        3401 => 8X"00",
        3402 => 8X"00",
        3403 => 8X"00",
        3404 => 8X"00",
        3405 => 8X"00",
        3406 => 8X"00",
        3407 => 8X"00",
        3408 => 8X"00",
        3409 => 8X"00",
        3410 => 8X"00",
        3411 => 8X"00",
        3412 => 8X"00",
        3413 => 8X"00",
        3414 => 8X"1F",
        3415 => 8X"18",
        3416 => 8X"1F",
        3417 => 8X"18",
        3418 => 8X"18",
        3419 => 8X"18",
        3420 => 8X"18",
        3421 => 8X"18",
        3422 => 8X"18",
        3423 => 8X"18",
        3424 => 8X"00",
        3425 => 8X"00",
        3426 => 8X"00",
        3427 => 8X"00",
        3428 => 8X"00",
        3429 => 8X"00",
        3430 => 8X"00",
        3431 => 8X"00",
        3432 => 8X"3F",
        3433 => 8X"36",
        3434 => 8X"36",
        3435 => 8X"36",
        3436 => 8X"36",
        3437 => 8X"36",
        3438 => 8X"36",
        3439 => 8X"36",
        3440 => 8X"36",
        3441 => 8X"36",
        3442 => 8X"36",
        3443 => 8X"36",
        3444 => 8X"36",
        3445 => 8X"36",
        3446 => 8X"36",
        3447 => 8X"36",
        3448 => 8X"FF",
        3449 => 8X"36",
        3450 => 8X"36",
        3451 => 8X"36",
        3452 => 8X"36",
        3453 => 8X"36",
        3454 => 8X"36",
        3455 => 8X"36",
        3456 => 8X"18",
        3457 => 8X"18",
        3458 => 8X"18",
        3459 => 8X"18",
        3460 => 8X"18",
        3461 => 8X"18",
        3462 => 8X"FF",
        3463 => 8X"18",
        3464 => 8X"FF",
        3465 => 8X"18",
        3466 => 8X"18",
        3467 => 8X"18",
        3468 => 8X"18",
        3469 => 8X"18",
        3470 => 8X"18",
        3471 => 8X"18",
        3472 => 8X"18",
        3473 => 8X"18",
        3474 => 8X"18",
        3475 => 8X"18",
        3476 => 8X"18",
        3477 => 8X"18",
        3478 => 8X"18",
        3479 => 8X"18",
        3480 => 8X"F8",
        3481 => 8X"00",
        3482 => 8X"00",
        3483 => 8X"00",
        3484 => 8X"00",
        3485 => 8X"00",
        3486 => 8X"00",
        3487 => 8X"00",
        3488 => 8X"00",
        3489 => 8X"00",
        3490 => 8X"00",
        3491 => 8X"00",
        3492 => 8X"00",
        3493 => 8X"00",
        3494 => 8X"00",
        3495 => 8X"00",
        3496 => 8X"1F",
        3497 => 8X"18",
        3498 => 8X"18",
        3499 => 8X"18",
        3500 => 8X"18",
        3501 => 8X"18",
        3502 => 8X"18",
        3503 => 8X"18",
        3504 => 8X"FF",
        3505 => 8X"FF",
        3506 => 8X"FF",
        3507 => 8X"FF",
        3508 => 8X"FF",
        3509 => 8X"FF",
        3510 => 8X"FF",
        3511 => 8X"FF",
        3512 => 8X"FF",
        3513 => 8X"FF",
        3514 => 8X"FF",
        3515 => 8X"FF",
        3516 => 8X"FF",
        3517 => 8X"FF",
        3518 => 8X"FF",
        3519 => 8X"FF",
        3520 => 8X"00",
        3521 => 8X"00",
        3522 => 8X"00",
        3523 => 8X"00",
        3524 => 8X"00",
        3525 => 8X"00",
        3526 => 8X"00",
        3527 => 8X"00",
        3528 => 8X"FF",
        3529 => 8X"FF",
        3530 => 8X"FF",
        3531 => 8X"FF",
        3532 => 8X"FF",
        3533 => 8X"FF",
        3534 => 8X"FF",
        3535 => 8X"FF",
        3536 => 8X"F0",
        3537 => 8X"F0",
        3538 => 8X"F0",
        3539 => 8X"F0",
        3540 => 8X"F0",
        3541 => 8X"F0",
        3542 => 8X"F0",
        3543 => 8X"F0",
        3544 => 8X"F0",
        3545 => 8X"F0",
        3546 => 8X"F0",
        3547 => 8X"F0",
        3548 => 8X"F0",
        3549 => 8X"F0",
        3550 => 8X"F0",
        3551 => 8X"F0",
        3552 => 8X"0F",
        3553 => 8X"0F",
        3554 => 8X"0F",
        3555 => 8X"0F",
        3556 => 8X"0F",
        3557 => 8X"0F",
        3558 => 8X"0F",
        3559 => 8X"0F",
        3560 => 8X"0F",
        3561 => 8X"0F",
        3562 => 8X"0F",
        3563 => 8X"0F",
        3564 => 8X"0F",
        3565 => 8X"0F",
        3566 => 8X"0F",
        3567 => 8X"0F",
        3568 => 8X"FF",
        3569 => 8X"FF",
        3570 => 8X"FF",
        3571 => 8X"FF",
        3572 => 8X"FF",
        3573 => 8X"FF",
        3574 => 8X"FF",
        3575 => 8X"FF",
        3576 => 8X"00",
        3577 => 8X"00",
        3578 => 8X"00",
        3579 => 8X"00",
        3580 => 8X"00",
        3581 => 8X"00",
        3582 => 8X"00",
        3583 => 8X"00",
        3584 => 8X"00",
        3585 => 8X"00",
        3586 => 8X"00",
        3587 => 8X"00",
        3588 => 8X"00",
        3589 => 8X"DC",
        3590 => 8X"66",
        3591 => 8X"66",
        3592 => 8X"66",
        3593 => 8X"66",
        3594 => 8X"66",
        3595 => 8X"7C",
        3596 => 8X"60",
        3597 => 8X"60",
        3598 => 8X"F0",
        3599 => 8X"00",
        3600 => 8X"00",
        3601 => 8X"00",
        3602 => 8X"00",
        3603 => 8X"00",
        3604 => 8X"00",
        3605 => 8X"7C",
        3606 => 8X"C6",
        3607 => 8X"C6",
        3608 => 8X"C0",
        3609 => 8X"C0",
        3610 => 8X"C6",
        3611 => 8X"C6",
        3612 => 8X"7C",
        3613 => 8X"00",
        3614 => 8X"00",
        3615 => 8X"00",
        3616 => 8X"00",
        3617 => 8X"00",
        3618 => 8X"00",
        3619 => 8X"00",
        3620 => 8X"00",
        3621 => 8X"7E",
        3622 => 8X"5A",
        3623 => 8X"18",
        3624 => 8X"18",
        3625 => 8X"18",
        3626 => 8X"18",
        3627 => 8X"18",
        3628 => 8X"3C",
        3629 => 8X"00",
        3630 => 8X"00",
        3631 => 8X"00",
        3632 => 8X"00",
        3633 => 8X"00",
        3634 => 8X"00",
        3635 => 8X"00",
        3636 => 8X"00",
        3637 => 8X"C6",
        3638 => 8X"C6",
        3639 => 8X"C6",
        3640 => 8X"C6",
        3641 => 8X"C6",
        3642 => 8X"C6",
        3643 => 8X"7E",
        3644 => 8X"06",
        3645 => 8X"0C",
        3646 => 8X"F8",
        3647 => 8X"00",
        3648 => 8X"00",
        3649 => 8X"00",
        3650 => 8X"00",
        3651 => 8X"00",
        3652 => 8X"00",
        3653 => 8X"18",
        3654 => 8X"7E",
        3655 => 8X"DB",
        3656 => 8X"DB",
        3657 => 8X"DB",
        3658 => 8X"DB",
        3659 => 8X"DB",
        3660 => 8X"7E",
        3661 => 8X"18",
        3662 => 8X"18",
        3663 => 8X"00",
        3664 => 8X"00",
        3665 => 8X"00",
        3666 => 8X"00",
        3667 => 8X"00",
        3668 => 8X"00",
        3669 => 8X"C6",
        3670 => 8X"C6",
        3671 => 8X"6C",
        3672 => 8X"38",
        3673 => 8X"38",
        3674 => 8X"6C",
        3675 => 8X"C6",
        3676 => 8X"C6",
        3677 => 8X"00",
        3678 => 8X"00",
        3679 => 8X"00",
        3680 => 8X"00",
        3681 => 8X"00",
        3682 => 8X"00",
        3683 => 8X"00",
        3684 => 8X"00",
        3685 => 8X"CC",
        3686 => 8X"CC",
        3687 => 8X"CC",
        3688 => 8X"CC",
        3689 => 8X"CC",
        3690 => 8X"CC",
        3691 => 8X"CC",
        3692 => 8X"FE",
        3693 => 8X"06",
        3694 => 8X"06",
        3695 => 8X"00",
        3696 => 8X"00",
        3697 => 8X"00",
        3698 => 8X"00",
        3699 => 8X"00",
        3700 => 8X"00",
        3701 => 8X"C6",
        3702 => 8X"C6",
        3703 => 8X"C6",
        3704 => 8X"C6",
        3705 => 8X"7E",
        3706 => 8X"06",
        3707 => 8X"06",
        3708 => 8X"06",
        3709 => 8X"00",
        3710 => 8X"00",
        3711 => 8X"00",
        3712 => 8X"00",
        3713 => 8X"00",
        3714 => 8X"00",
        3715 => 8X"00",
        3716 => 8X"00",
        3717 => 8X"D6",
        3718 => 8X"D6",
        3719 => 8X"D6",
        3720 => 8X"D6",
        3721 => 8X"D6",
        3722 => 8X"D6",
        3723 => 8X"D6",
        3724 => 8X"FE",
        3725 => 8X"00",
        3726 => 8X"00",
        3727 => 8X"00",
        3728 => 8X"00",
        3729 => 8X"00",
        3730 => 8X"00",
        3731 => 8X"00",
        3732 => 8X"00",
        3733 => 8X"D6",
        3734 => 8X"D6",
        3735 => 8X"D6",
        3736 => 8X"D6",
        3737 => 8X"D6",
        3738 => 8X"D6",
        3739 => 8X"D6",
        3740 => 8X"FE",
        3741 => 8X"03",
        3742 => 8X"03",
        3743 => 8X"00",
        3744 => 8X"00",
        3745 => 8X"00",
        3746 => 8X"00",
        3747 => 8X"00",
        3748 => 8X"00",
        3749 => 8X"F8",
        3750 => 8X"B0",
        3751 => 8X"3C",
        3752 => 8X"36",
        3753 => 8X"36",
        3754 => 8X"36",
        3755 => 8X"36",
        3756 => 8X"7C",
        3757 => 8X"00",
        3758 => 8X"00",
        3759 => 8X"00",
        3760 => 8X"00",
        3761 => 8X"00",
        3762 => 8X"00",
        3763 => 8X"00",
        3764 => 8X"00",
        3765 => 8X"C6",
        3766 => 8X"C6",
        3767 => 8X"F6",
        3768 => 8X"DE",
        3769 => 8X"DE",
        3770 => 8X"DE",
        3771 => 8X"DE",
        3772 => 8X"F6",
        3773 => 8X"00",
        3774 => 8X"00",
        3775 => 8X"00",
        3776 => 8X"00",
        3777 => 8X"00",
        3778 => 8X"00",
        3779 => 8X"00",
        3780 => 8X"00",
        3781 => 8X"F0",
        3782 => 8X"60",
        3783 => 8X"60",
        3784 => 8X"7C",
        3785 => 8X"66",
        3786 => 8X"66",
        3787 => 8X"66",
        3788 => 8X"FC",
        3789 => 8X"00",
        3790 => 8X"00",
        3791 => 8X"00",
        3792 => 8X"00",
        3793 => 8X"00",
        3794 => 8X"00",
        3795 => 8X"00",
        3796 => 8X"00",
        3797 => 8X"3C",
        3798 => 8X"66",
        3799 => 8X"06",
        3800 => 8X"1E",
        3801 => 8X"06",
        3802 => 8X"66",
        3803 => 8X"66",
        3804 => 8X"3C",
        3805 => 8X"00",
        3806 => 8X"00",
        3807 => 8X"00",
        3808 => 8X"00",
        3809 => 8X"00",
        3810 => 8X"00",
        3811 => 8X"00",
        3812 => 8X"00",
        3813 => 8X"9C",
        3814 => 8X"B6",
        3815 => 8X"B6",
        3816 => 8X"F6",
        3817 => 8X"B6",
        3818 => 8X"B6",
        3819 => 8X"B6",
        3820 => 8X"9C",
        3821 => 8X"00",
        3822 => 8X"00",
        3823 => 8X"00",
        3824 => 8X"00",
        3825 => 8X"00",
        3826 => 8X"00",
        3827 => 8X"00",
        3828 => 8X"00",
        3829 => 8X"7E",
        3830 => 8X"CC",
        3831 => 8X"CC",
        3832 => 8X"CC",
        3833 => 8X"7C",
        3834 => 8X"6C",
        3835 => 8X"CC",
        3836 => 8X"CE",
        3837 => 8X"00",
        3838 => 8X"00",
        3839 => 8X"00",
        3840 => 8X"00",
        3841 => 8X"00",
        3842 => 8X"00",
        3843 => 8X"00",
        3844 => 8X"FE",
        3845 => 8X"00",
        3846 => 8X"00",
        3847 => 8X"FE",
        3848 => 8X"00",
        3849 => 8X"00",
        3850 => 8X"FE",
        3851 => 8X"00",
        3852 => 8X"00",
        3853 => 8X"00",
        3854 => 8X"00",
        3855 => 8X"00",
        3856 => 8X"00",
        3857 => 8X"00",
        3858 => 8X"00",
        3859 => 8X"00",
        3860 => 8X"18",
        3861 => 8X"18",
        3862 => 8X"7E",
        3863 => 8X"18",
        3864 => 8X"18",
        3865 => 8X"00",
        3866 => 8X"00",
        3867 => 8X"FF",
        3868 => 8X"00",
        3869 => 8X"00",
        3870 => 8X"00",
        3871 => 8X"00",
        3872 => 8X"00",
        3873 => 8X"00",
        3874 => 8X"00",
        3875 => 8X"30",
        3876 => 8X"18",
        3877 => 8X"0C",
        3878 => 8X"06",
        3879 => 8X"0C",
        3880 => 8X"18",
        3881 => 8X"30",
        3882 => 8X"00",
        3883 => 8X"7E",
        3884 => 8X"00",
        3885 => 8X"00",
        3886 => 8X"00",
        3887 => 8X"00",
        3888 => 8X"00",
        3889 => 8X"00",
        3890 => 8X"00",
        3891 => 8X"0C",
        3892 => 8X"18",
        3893 => 8X"30",
        3894 => 8X"60",
        3895 => 8X"30",
        3896 => 8X"18",
        3897 => 8X"0C",
        3898 => 8X"00",
        3899 => 8X"7E",
        3900 => 8X"00",
        3901 => 8X"00",
        3902 => 8X"00",
        3903 => 8X"00",
        3904 => 8X"00",
        3905 => 8X"00",
        3906 => 8X"00",
        3907 => 8X"0E",
        3908 => 8X"1B",
        3909 => 8X"1B",
        3910 => 8X"18",
        3911 => 8X"18",
        3912 => 8X"18",
        3913 => 8X"18",
        3914 => 8X"18",
        3915 => 8X"18",
        3916 => 8X"18",
        3917 => 8X"18",
        3918 => 8X"18",
        3919 => 8X"18",
        3920 => 8X"18",
        3921 => 8X"18",
        3922 => 8X"18",
        3923 => 8X"18",
        3924 => 8X"18",
        3925 => 8X"18",
        3926 => 8X"18",
        3927 => 8X"18",
        3928 => 8X"18",
        3929 => 8X"D8",
        3930 => 8X"D8",
        3931 => 8X"70",
        3932 => 8X"00",
        3933 => 8X"00",
        3934 => 8X"00",
        3935 => 8X"00",
        3936 => 8X"00",
        3937 => 8X"00",
        3938 => 8X"00",
        3939 => 8X"00",
        3940 => 8X"18",
        3941 => 8X"18",
        3942 => 8X"00",
        3943 => 8X"7E",
        3944 => 8X"00",
        3945 => 8X"18",
        3946 => 8X"18",
        3947 => 8X"00",
        3948 => 8X"00",
        3949 => 8X"00",
        3950 => 8X"00",
        3951 => 8X"00",
        3952 => 8X"00",
        3953 => 8X"00",
        3954 => 8X"00",
        3955 => 8X"00",
        3956 => 8X"00",
        3957 => 8X"76",
        3958 => 8X"DC",
        3959 => 8X"00",
        3960 => 8X"76",
        3961 => 8X"DC",
        3962 => 8X"00",
        3963 => 8X"00",
        3964 => 8X"00",
        3965 => 8X"00",
        3966 => 8X"00",
        3967 => 8X"00",
        3968 => 8X"00",
        3969 => 8X"38",
        3970 => 8X"6C",
        3971 => 8X"6C",
        3972 => 8X"6C",
        3973 => 8X"38",
        3974 => 8X"00",
        3975 => 8X"00",
        3976 => 8X"00",
        3977 => 8X"00",
        3978 => 8X"00",
        3979 => 8X"00",
        3980 => 8X"00",
        3981 => 8X"00",
        3982 => 8X"00",
        3983 => 8X"00",
        3984 => 8X"00",
        3985 => 8X"00",
        3986 => 8X"00",
        3987 => 8X"00",
        3988 => 8X"00",
        3989 => 8X"00",
        3990 => 8X"00",
        3991 => 8X"18",
        3992 => 8X"18",
        3993 => 8X"00",
        3994 => 8X"00",
        3995 => 8X"00",
        3996 => 8X"00",
        3997 => 8X"00",
        3998 => 8X"00",
        3999 => 8X"00",
        4000 => 8X"00",
        4001 => 8X"00",
        4002 => 8X"00",
        4003 => 8X"00",
        4004 => 8X"00",
        4005 => 8X"00",
        4006 => 8X"00",
        4007 => 8X"00",
        4008 => 8X"18",
        4009 => 8X"00",
        4010 => 8X"00",
        4011 => 8X"00",
        4012 => 8X"00",
        4013 => 8X"00",
        4014 => 8X"00",
        4015 => 8X"00",
        4016 => 8X"00",
        4017 => 8X"0F",
        4018 => 8X"0C",
        4019 => 8X"0C",
        4020 => 8X"0C",
        4021 => 8X"0C",
        4022 => 8X"0C",
        4023 => 8X"EC",
        4024 => 8X"6C",
        4025 => 8X"3C",
        4026 => 8X"1C",
        4027 => 8X"0C",
        4028 => 8X"00",
        4029 => 8X"00",
        4030 => 8X"00",
        4031 => 8X"00",
        4032 => 8X"00",
        4033 => 8X"00",
        4034 => 8X"D8",
        4035 => 8X"6C",
        4036 => 8X"6C",
        4037 => 8X"6C",
        4038 => 8X"6C",
        4039 => 8X"6C",
        4040 => 8X"00",
        4041 => 8X"00",
        4042 => 8X"00",
        4043 => 8X"00",
        4044 => 8X"00",
        4045 => 8X"00",
        4046 => 8X"00",
        4047 => 8X"00",
        4048 => 8X"00",
        4049 => 8X"00",
        4050 => 8X"70",
        4051 => 8X"D8",
        4052 => 8X"30",
        4053 => 8X"60",
        4054 => 8X"C8",
        4055 => 8X"F8",
        4056 => 8X"00",
        4057 => 8X"00",
        4058 => 8X"00",
        4059 => 8X"00",
        4060 => 8X"00",
        4061 => 8X"00",
        4062 => 8X"00",
        4063 => 8X"00",
        4064 => 8X"00",
        4065 => 8X"00",
        4066 => 8X"00",
        4067 => 8X"00",
        4068 => 8X"3C",
        4069 => 8X"3C",
        4070 => 8X"3C",
        4071 => 8X"3C",
        4072 => 8X"3C",
        4073 => 8X"3C",
        4074 => 8X"3C",
        4075 => 8X"3C",
        4076 => 8X"00",
        4077 => 8X"00",
        4078 => 8X"00",
        4079 => 8X"00",
        4080 => 8X"00",
        4081 => 8X"00",
        4082 => 8X"00",
        4083 => 8X"00",
        4084 => 8X"00",
        4085 => 8X"00",
        4086 => 8X"00",
        4087 => 8X"00",
        4088 => 8X"00",
        4089 => 8X"00",
        4090 => 8X"00",
        4091 => 8X"00",
        4092 => 8X"00",
        4093 => 8X"00",
        4094 => 8X"00",
        4095 => 8X"00",
        others => X"XX"
    );

end package symbol_mem_pkg;
