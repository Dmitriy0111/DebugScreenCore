--
-- File            :   display_mem_schoolMIPS_pkg.vhd
-- Autor           :   Vlasov D.V.
-- Data            :   2019.06.10
-- Language        :   VHDL
-- Description     :   This display memory file for DebugScreenCore for schoolMIPS
-- Copyright(c)    :   2019 Vlasov D.V.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library dsc;
use dsc.dsc_mem_pkg.all;

package display_mem_schoolMIPS_pkg is

    constant display_mem_schoolMIPS_hex : mem_t(2559 downto 0)(7 downto 0) :=
    (
           0 => 8X"70",
           1 => 8X"63",
           2 => 8X"3A",
           3 => 8X"20",
           4 => 8X"30",
           5 => 8X"78",
           6 => 8X"2A",
           7 => 8X"2A",
           8 => 8X"2A",
           9 => 8X"2A",
          10 => 8X"2A",
          11 => 8X"2A",
          12 => 8X"2A",
          13 => 8X"2A",
          14 => 8X"20",
          15 => 8X"20",
          16 => 8X"20",
          17 => 8X"20",
          18 => 8X"20",
          19 => 8X"20",
          20 => 8X"20",
          21 => 8X"20",
          22 => 8X"20",
          23 => 8X"20",
          24 => 8X"20",
          25 => 8X"20",
          26 => 8X"20",
          27 => 8X"20",
          28 => 8X"20",
          29 => 8X"20",
          30 => 8X"20",
          31 => 8X"20",
          32 => 8X"20",
          33 => 8X"20",
          34 => 8X"20",
          35 => 8X"20",
          36 => 8X"20",
          37 => 8X"20",
          38 => 8X"20",
          39 => 8X"20",
          40 => 8X"20",
          41 => 8X"20",
          42 => 8X"20",
          43 => 8X"20",
          44 => 8X"20",
          45 => 8X"20",
          46 => 8X"20",
          47 => 8X"20",
          48 => 8X"20",
          49 => 8X"20",
          50 => 8X"20",
          51 => 8X"20",
          52 => 8X"54",
          53 => 8X"68",
          54 => 8X"69",
          55 => 8X"73",
          56 => 8X"20",
          57 => 8X"69",
          58 => 8X"73",
          59 => 8X"20",
          60 => 8X"53",
          61 => 8X"63",
          62 => 8X"68",
          63 => 8X"6F",
          64 => 8X"6F",
          65 => 8X"6C",
          66 => 8X"4D",
          67 => 8X"49",
          68 => 8X"50",
          69 => 8X"53",
          70 => 8X"20",
          71 => 8X"72",
          72 => 8X"65",
          73 => 8X"67",
          74 => 8X"69",
          75 => 8X"73",
          76 => 8X"74",
          77 => 8X"65",
          78 => 8X"72",
          79 => 8X"73",
          80 => 8X"61",
          81 => 8X"74",
          82 => 8X"3A",
          83 => 8X"20",
          84 => 8X"30",
          85 => 8X"78",
          86 => 8X"2A",
          87 => 8X"2A",
          88 => 8X"2A",
          89 => 8X"2A",
          90 => 8X"2A",
          91 => 8X"2A",
          92 => 8X"2A",
          93 => 8X"2A",
          94 => 8X"20",
          95 => 8X"20",
          96 => 8X"20",
          97 => 8X"20",
          98 => 8X"20",
          99 => 8X"20",
         100 => 8X"20",
         101 => 8X"20",
         102 => 8X"20",
         103 => 8X"20",
         104 => 8X"20",
         105 => 8X"20",
         106 => 8X"20",
         107 => 8X"20",
         108 => 8X"20",
         109 => 8X"20",
         110 => 8X"20",
         111 => 8X"20",
         112 => 8X"20",
         113 => 8X"20",
         114 => 8X"20",
         115 => 8X"20",
         116 => 8X"20",
         117 => 8X"20",
         118 => 8X"20",
         119 => 8X"20",
         120 => 8X"20",
         121 => 8X"20",
         122 => 8X"20",
         123 => 8X"20",
         124 => 8X"20",
         125 => 8X"20",
         126 => 8X"20",
         127 => 8X"20",
         128 => 8X"20",
         129 => 8X"20",
         130 => 8X"20",
         131 => 8X"20",
         132 => 8X"20",
         133 => 8X"20",
         134 => 8X"20",
         135 => 8X"20",
         136 => 8X"20",
         137 => 8X"20",
         138 => 8X"20",
         139 => 8X"20",
         140 => 8X"20",
         141 => 8X"20",
         142 => 8X"20",
         143 => 8X"20",
         144 => 8X"20",
         145 => 8X"20",
         146 => 8X"20",
         147 => 8X"20",
         148 => 8X"20",
         149 => 8X"20",
         150 => 8X"20",
         151 => 8X"20",
         152 => 8X"20",
         153 => 8X"20",
         154 => 8X"20",
         155 => 8X"20",
         156 => 8X"20",
         157 => 8X"20",
         158 => 8X"20",
         159 => 8X"20",
         160 => 8X"76",
         161 => 8X"30",
         162 => 8X"3A",
         163 => 8X"20",
         164 => 8X"30",
         165 => 8X"78",
         166 => 8X"2A",
         167 => 8X"2A",
         168 => 8X"2A",
         169 => 8X"2A",
         170 => 8X"2A",
         171 => 8X"2A",
         172 => 8X"2A",
         173 => 8X"2A",
         174 => 8X"20",
         175 => 8X"20",
         176 => 8X"20",
         177 => 8X"20",
         178 => 8X"20",
         179 => 8X"20",
         180 => 8X"20",
         181 => 8X"20",
         182 => 8X"20",
         183 => 8X"20",
         184 => 8X"20",
         185 => 8X"20",
         186 => 8X"20",
         187 => 8X"20",
         188 => 8X"20",
         189 => 8X"20",
         190 => 8X"20",
         191 => 8X"20",
         192 => 8X"20",
         193 => 8X"20",
         194 => 8X"20",
         195 => 8X"20",
         196 => 8X"20",
         197 => 8X"20",
         198 => 8X"20",
         199 => 8X"20",
         200 => 8X"20",
         201 => 8X"20",
         202 => 8X"20",
         203 => 8X"20",
         204 => 8X"20",
         205 => 8X"20",
         206 => 8X"20",
         207 => 8X"20",
         208 => 8X"20",
         209 => 8X"20",
         210 => 8X"20",
         211 => 8X"20",
         212 => 8X"20",
         213 => 8X"20",
         214 => 8X"20",
         215 => 8X"20",
         216 => 8X"20",
         217 => 8X"20",
         218 => 8X"20",
         219 => 8X"20",
         220 => 8X"20",
         221 => 8X"20",
         222 => 8X"20",
         223 => 8X"20",
         224 => 8X"20",
         225 => 8X"20",
         226 => 8X"20",
         227 => 8X"20",
         228 => 8X"20",
         229 => 8X"20",
         230 => 8X"20",
         231 => 8X"20",
         232 => 8X"20",
         233 => 8X"20",
         234 => 8X"20",
         235 => 8X"20",
         236 => 8X"20",
         237 => 8X"20",
         238 => 8X"20",
         239 => 8X"20",
         240 => 8X"76",
         241 => 8X"31",
         242 => 8X"3A",
         243 => 8X"20",
         244 => 8X"30",
         245 => 8X"78",
         246 => 8X"2A",
         247 => 8X"2A",
         248 => 8X"2A",
         249 => 8X"2A",
         250 => 8X"2A",
         251 => 8X"2A",
         252 => 8X"2A",
         253 => 8X"2A",
         254 => 8X"20",
         255 => 8X"20",
         256 => 8X"20",
         257 => 8X"20",
         258 => 8X"20",
         259 => 8X"20",
         260 => 8X"20",
         261 => 8X"20",
         262 => 8X"20",
         263 => 8X"20",
         264 => 8X"20",
         265 => 8X"20",
         266 => 8X"20",
         267 => 8X"20",
         268 => 8X"20",
         269 => 8X"20",
         270 => 8X"20",
         271 => 8X"20",
         272 => 8X"20",
         273 => 8X"20",
         274 => 8X"20",
         275 => 8X"20",
         276 => 8X"20",
         277 => 8X"20",
         278 => 8X"20",
         279 => 8X"20",
         280 => 8X"20",
         281 => 8X"20",
         282 => 8X"20",
         283 => 8X"20",
         284 => 8X"20",
         285 => 8X"20",
         286 => 8X"20",
         287 => 8X"20",
         288 => 8X"20",
         289 => 8X"20",
         290 => 8X"20",
         291 => 8X"20",
         292 => 8X"20",
         293 => 8X"20",
         294 => 8X"20",
         295 => 8X"20",
         296 => 8X"20",
         297 => 8X"20",
         298 => 8X"20",
         299 => 8X"20",
         300 => 8X"20",
         301 => 8X"20",
         302 => 8X"20",
         303 => 8X"20",
         304 => 8X"20",
         305 => 8X"20",
         306 => 8X"20",
         307 => 8X"20",
         308 => 8X"20",
         309 => 8X"20",
         310 => 8X"20",
         311 => 8X"20",
         312 => 8X"20",
         313 => 8X"20",
         314 => 8X"20",
         315 => 8X"20",
         316 => 8X"20",
         317 => 8X"20",
         318 => 8X"20",
         319 => 8X"20",
         320 => 8X"61",
         321 => 8X"30",
         322 => 8X"3A",
         323 => 8X"20",
         324 => 8X"30",
         325 => 8X"78",
         326 => 8X"2A",
         327 => 8X"2A",
         328 => 8X"2A",
         329 => 8X"2A",
         330 => 8X"2A",
         331 => 8X"2A",
         332 => 8X"2A",
         333 => 8X"2A",
         334 => 8X"20",
         335 => 8X"20",
         336 => 8X"20",
         337 => 8X"20",
         338 => 8X"20",
         339 => 8X"20",
         340 => 8X"20",
         341 => 8X"20",
         342 => 8X"20",
         343 => 8X"20",
         344 => 8X"20",
         345 => 8X"20",
         346 => 8X"20",
         347 => 8X"20",
         348 => 8X"20",
         349 => 8X"20",
         350 => 8X"20",
         351 => 8X"20",
         352 => 8X"20",
         353 => 8X"20",
         354 => 8X"20",
         355 => 8X"20",
         356 => 8X"20",
         357 => 8X"20",
         358 => 8X"20",
         359 => 8X"20",
         360 => 8X"20",
         361 => 8X"20",
         362 => 8X"20",
         363 => 8X"20",
         364 => 8X"20",
         365 => 8X"20",
         366 => 8X"20",
         367 => 8X"20",
         368 => 8X"20",
         369 => 8X"20",
         370 => 8X"20",
         371 => 8X"20",
         372 => 8X"20",
         373 => 8X"20",
         374 => 8X"20",
         375 => 8X"20",
         376 => 8X"20",
         377 => 8X"20",
         378 => 8X"20",
         379 => 8X"20",
         380 => 8X"20",
         381 => 8X"20",
         382 => 8X"20",
         383 => 8X"20",
         384 => 8X"20",
         385 => 8X"20",
         386 => 8X"20",
         387 => 8X"20",
         388 => 8X"20",
         389 => 8X"20",
         390 => 8X"20",
         391 => 8X"20",
         392 => 8X"20",
         393 => 8X"20",
         394 => 8X"20",
         395 => 8X"20",
         396 => 8X"20",
         397 => 8X"20",
         398 => 8X"20",
         399 => 8X"20",
         400 => 8X"61",
         401 => 8X"31",
         402 => 8X"3A",
         403 => 8X"20",
         404 => 8X"30",
         405 => 8X"78",
         406 => 8X"2A",
         407 => 8X"2A",
         408 => 8X"2A",
         409 => 8X"2A",
         410 => 8X"2A",
         411 => 8X"2A",
         412 => 8X"2A",
         413 => 8X"2A",
         414 => 8X"20",
         415 => 8X"20",
         416 => 8X"20",
         417 => 8X"20",
         418 => 8X"20",
         419 => 8X"20",
         420 => 8X"20",
         421 => 8X"20",
         422 => 8X"20",
         423 => 8X"20",
         424 => 8X"20",
         425 => 8X"20",
         426 => 8X"20",
         427 => 8X"20",
         428 => 8X"20",
         429 => 8X"20",
         430 => 8X"20",
         431 => 8X"20",
         432 => 8X"20",
         433 => 8X"20",
         434 => 8X"20",
         435 => 8X"20",
         436 => 8X"20",
         437 => 8X"20",
         438 => 8X"20",
         439 => 8X"20",
         440 => 8X"20",
         441 => 8X"20",
         442 => 8X"20",
         443 => 8X"20",
         444 => 8X"20",
         445 => 8X"20",
         446 => 8X"20",
         447 => 8X"20",
         448 => 8X"20",
         449 => 8X"20",
         450 => 8X"20",
         451 => 8X"20",
         452 => 8X"20",
         453 => 8X"20",
         454 => 8X"20",
         455 => 8X"20",
         456 => 8X"20",
         457 => 8X"20",
         458 => 8X"20",
         459 => 8X"20",
         460 => 8X"20",
         461 => 8X"20",
         462 => 8X"20",
         463 => 8X"20",
         464 => 8X"20",
         465 => 8X"20",
         466 => 8X"20",
         467 => 8X"20",
         468 => 8X"20",
         469 => 8X"20",
         470 => 8X"20",
         471 => 8X"20",
         472 => 8X"20",
         473 => 8X"20",
         474 => 8X"20",
         475 => 8X"20",
         476 => 8X"20",
         477 => 8X"20",
         478 => 8X"20",
         479 => 8X"20",
         480 => 8X"61",
         481 => 8X"32",
         482 => 8X"3A",
         483 => 8X"20",
         484 => 8X"30",
         485 => 8X"78",
         486 => 8X"2A",
         487 => 8X"2A",
         488 => 8X"2A",
         489 => 8X"2A",
         490 => 8X"2A",
         491 => 8X"2A",
         492 => 8X"2A",
         493 => 8X"2A",
         494 => 8X"20",
         495 => 8X"20",
         496 => 8X"20",
         497 => 8X"20",
         498 => 8X"20",
         499 => 8X"20",
         500 => 8X"20",
         501 => 8X"20",
         502 => 8X"20",
         503 => 8X"20",
         504 => 8X"20",
         505 => 8X"20",
         506 => 8X"20",
         507 => 8X"20",
         508 => 8X"20",
         509 => 8X"20",
         510 => 8X"20",
         511 => 8X"20",
         512 => 8X"20",
         513 => 8X"20",
         514 => 8X"20",
         515 => 8X"20",
         516 => 8X"20",
         517 => 8X"20",
         518 => 8X"20",
         519 => 8X"20",
         520 => 8X"20",
         521 => 8X"20",
         522 => 8X"20",
         523 => 8X"20",
         524 => 8X"20",
         525 => 8X"20",
         526 => 8X"20",
         527 => 8X"20",
         528 => 8X"20",
         529 => 8X"20",
         530 => 8X"20",
         531 => 8X"20",
         532 => 8X"20",
         533 => 8X"20",
         534 => 8X"20",
         535 => 8X"20",
         536 => 8X"20",
         537 => 8X"20",
         538 => 8X"20",
         539 => 8X"20",
         540 => 8X"20",
         541 => 8X"20",
         542 => 8X"20",
         543 => 8X"20",
         544 => 8X"20",
         545 => 8X"20",
         546 => 8X"20",
         547 => 8X"20",
         548 => 8X"20",
         549 => 8X"20",
         550 => 8X"20",
         551 => 8X"20",
         552 => 8X"20",
         553 => 8X"20",
         554 => 8X"20",
         555 => 8X"20",
         556 => 8X"20",
         557 => 8X"20",
         558 => 8X"20",
         559 => 8X"20",
         560 => 8X"61",
         561 => 8X"33",
         562 => 8X"3A",
         563 => 8X"20",
         564 => 8X"30",
         565 => 8X"78",
         566 => 8X"2A",
         567 => 8X"2A",
         568 => 8X"2A",
         569 => 8X"2A",
         570 => 8X"2A",
         571 => 8X"2A",
         572 => 8X"2A",
         573 => 8X"2A",
         574 => 8X"20",
         575 => 8X"20",
         576 => 8X"20",
         577 => 8X"20",
         578 => 8X"20",
         579 => 8X"20",
         580 => 8X"20",
         581 => 8X"20",
         582 => 8X"20",
         583 => 8X"20",
         584 => 8X"20",
         585 => 8X"20",
         586 => 8X"20",
         587 => 8X"20",
         588 => 8X"20",
         589 => 8X"20",
         590 => 8X"20",
         591 => 8X"20",
         592 => 8X"20",
         593 => 8X"20",
         594 => 8X"20",
         595 => 8X"20",
         596 => 8X"20",
         597 => 8X"20",
         598 => 8X"20",
         599 => 8X"20",
         600 => 8X"20",
         601 => 8X"20",
         602 => 8X"20",
         603 => 8X"20",
         604 => 8X"20",
         605 => 8X"20",
         606 => 8X"20",
         607 => 8X"20",
         608 => 8X"20",
         609 => 8X"20",
         610 => 8X"20",
         611 => 8X"20",
         612 => 8X"20",
         613 => 8X"20",
         614 => 8X"20",
         615 => 8X"20",
         616 => 8X"20",
         617 => 8X"20",
         618 => 8X"20",
         619 => 8X"20",
         620 => 8X"20",
         621 => 8X"20",
         622 => 8X"20",
         623 => 8X"20",
         624 => 8X"20",
         625 => 8X"20",
         626 => 8X"20",
         627 => 8X"20",
         628 => 8X"20",
         629 => 8X"20",
         630 => 8X"20",
         631 => 8X"20",
         632 => 8X"20",
         633 => 8X"20",
         634 => 8X"20",
         635 => 8X"20",
         636 => 8X"20",
         637 => 8X"20",
         638 => 8X"20",
         639 => 8X"20",
         640 => 8X"74",
         641 => 8X"30",
         642 => 8X"3A",
         643 => 8X"20",
         644 => 8X"30",
         645 => 8X"78",
         646 => 8X"2A",
         647 => 8X"2A",
         648 => 8X"2A",
         649 => 8X"2A",
         650 => 8X"2A",
         651 => 8X"2A",
         652 => 8X"2A",
         653 => 8X"2A",
         654 => 8X"20",
         655 => 8X"20",
         656 => 8X"20",
         657 => 8X"20",
         658 => 8X"20",
         659 => 8X"20",
         660 => 8X"20",
         661 => 8X"20",
         662 => 8X"20",
         663 => 8X"20",
         664 => 8X"20",
         665 => 8X"20",
         666 => 8X"20",
         667 => 8X"20",
         668 => 8X"20",
         669 => 8X"20",
         670 => 8X"20",
         671 => 8X"20",
         672 => 8X"20",
         673 => 8X"20",
         674 => 8X"20",
         675 => 8X"20",
         676 => 8X"20",
         677 => 8X"20",
         678 => 8X"20",
         679 => 8X"20",
         680 => 8X"20",
         681 => 8X"20",
         682 => 8X"20",
         683 => 8X"20",
         684 => 8X"20",
         685 => 8X"20",
         686 => 8X"20",
         687 => 8X"20",
         688 => 8X"20",
         689 => 8X"20",
         690 => 8X"20",
         691 => 8X"20",
         692 => 8X"20",
         693 => 8X"20",
         694 => 8X"20",
         695 => 8X"20",
         696 => 8X"20",
         697 => 8X"20",
         698 => 8X"20",
         699 => 8X"20",
         700 => 8X"20",
         701 => 8X"20",
         702 => 8X"20",
         703 => 8X"20",
         704 => 8X"20",
         705 => 8X"20",
         706 => 8X"20",
         707 => 8X"20",
         708 => 8X"20",
         709 => 8X"20",
         710 => 8X"20",
         711 => 8X"20",
         712 => 8X"20",
         713 => 8X"20",
         714 => 8X"20",
         715 => 8X"20",
         716 => 8X"20",
         717 => 8X"20",
         718 => 8X"20",
         719 => 8X"20",
         720 => 8X"74",
         721 => 8X"31",
         722 => 8X"3A",
         723 => 8X"20",
         724 => 8X"30",
         725 => 8X"78",
         726 => 8X"2A",
         727 => 8X"2A",
         728 => 8X"2A",
         729 => 8X"2A",
         730 => 8X"2A",
         731 => 8X"2A",
         732 => 8X"2A",
         733 => 8X"2A",
         734 => 8X"20",
         735 => 8X"20",
         736 => 8X"20",
         737 => 8X"20",
         738 => 8X"20",
         739 => 8X"20",
         740 => 8X"20",
         741 => 8X"20",
         742 => 8X"20",
         743 => 8X"20",
         744 => 8X"20",
         745 => 8X"20",
         746 => 8X"20",
         747 => 8X"20",
         748 => 8X"20",
         749 => 8X"20",
         750 => 8X"20",
         751 => 8X"20",
         752 => 8X"20",
         753 => 8X"20",
         754 => 8X"20",
         755 => 8X"20",
         756 => 8X"20",
         757 => 8X"20",
         758 => 8X"20",
         759 => 8X"20",
         760 => 8X"20",
         761 => 8X"20",
         762 => 8X"20",
         763 => 8X"20",
         764 => 8X"20",
         765 => 8X"20",
         766 => 8X"20",
         767 => 8X"20",
         768 => 8X"20",
         769 => 8X"20",
         770 => 8X"20",
         771 => 8X"20",
         772 => 8X"20",
         773 => 8X"20",
         774 => 8X"20",
         775 => 8X"20",
         776 => 8X"20",
         777 => 8X"20",
         778 => 8X"20",
         779 => 8X"20",
         780 => 8X"20",
         781 => 8X"20",
         782 => 8X"20",
         783 => 8X"20",
         784 => 8X"20",
         785 => 8X"20",
         786 => 8X"20",
         787 => 8X"20",
         788 => 8X"20",
         789 => 8X"20",
         790 => 8X"20",
         791 => 8X"20",
         792 => 8X"20",
         793 => 8X"20",
         794 => 8X"20",
         795 => 8X"20",
         796 => 8X"20",
         797 => 8X"20",
         798 => 8X"20",
         799 => 8X"20",
         800 => 8X"74",
         801 => 8X"32",
         802 => 8X"3A",
         803 => 8X"20",
         804 => 8X"30",
         805 => 8X"78",
         806 => 8X"2A",
         807 => 8X"2A",
         808 => 8X"2A",
         809 => 8X"2A",
         810 => 8X"2A",
         811 => 8X"2A",
         812 => 8X"2A",
         813 => 8X"2A",
         814 => 8X"20",
         815 => 8X"20",
         816 => 8X"20",
         817 => 8X"20",
         818 => 8X"20",
         819 => 8X"20",
         820 => 8X"20",
         821 => 8X"20",
         822 => 8X"20",
         823 => 8X"20",
         824 => 8X"20",
         825 => 8X"20",
         826 => 8X"20",
         827 => 8X"20",
         828 => 8X"20",
         829 => 8X"20",
         830 => 8X"20",
         831 => 8X"20",
         832 => 8X"20",
         833 => 8X"20",
         834 => 8X"20",
         835 => 8X"20",
         836 => 8X"20",
         837 => 8X"20",
         838 => 8X"20",
         839 => 8X"20",
         840 => 8X"20",
         841 => 8X"20",
         842 => 8X"20",
         843 => 8X"20",
         844 => 8X"20",
         845 => 8X"20",
         846 => 8X"20",
         847 => 8X"20",
         848 => 8X"20",
         849 => 8X"20",
         850 => 8X"20",
         851 => 8X"20",
         852 => 8X"20",
         853 => 8X"20",
         854 => 8X"20",
         855 => 8X"20",
         856 => 8X"20",
         857 => 8X"20",
         858 => 8X"20",
         859 => 8X"20",
         860 => 8X"20",
         861 => 8X"20",
         862 => 8X"20",
         863 => 8X"20",
         864 => 8X"20",
         865 => 8X"20",
         866 => 8X"20",
         867 => 8X"20",
         868 => 8X"20",
         869 => 8X"20",
         870 => 8X"20",
         871 => 8X"20",
         872 => 8X"20",
         873 => 8X"20",
         874 => 8X"20",
         875 => 8X"20",
         876 => 8X"20",
         877 => 8X"20",
         878 => 8X"20",
         879 => 8X"20",
         880 => 8X"74",
         881 => 8X"33",
         882 => 8X"3A",
         883 => 8X"20",
         884 => 8X"30",
         885 => 8X"78",
         886 => 8X"2A",
         887 => 8X"2A",
         888 => 8X"2A",
         889 => 8X"2A",
         890 => 8X"2A",
         891 => 8X"2A",
         892 => 8X"2A",
         893 => 8X"2A",
         894 => 8X"20",
         895 => 8X"20",
         896 => 8X"20",
         897 => 8X"20",
         898 => 8X"20",
         899 => 8X"20",
         900 => 8X"20",
         901 => 8X"20",
         902 => 8X"20",
         903 => 8X"20",
         904 => 8X"20",
         905 => 8X"20",
         906 => 8X"20",
         907 => 8X"20",
         908 => 8X"20",
         909 => 8X"20",
         910 => 8X"20",
         911 => 8X"20",
         912 => 8X"20",
         913 => 8X"20",
         914 => 8X"20",
         915 => 8X"20",
         916 => 8X"20",
         917 => 8X"20",
         918 => 8X"20",
         919 => 8X"20",
         920 => 8X"20",
         921 => 8X"20",
         922 => 8X"20",
         923 => 8X"20",
         924 => 8X"20",
         925 => 8X"20",
         926 => 8X"20",
         927 => 8X"20",
         928 => 8X"20",
         929 => 8X"20",
         930 => 8X"20",
         931 => 8X"20",
         932 => 8X"20",
         933 => 8X"20",
         934 => 8X"20",
         935 => 8X"20",
         936 => 8X"20",
         937 => 8X"20",
         938 => 8X"20",
         939 => 8X"20",
         940 => 8X"20",
         941 => 8X"20",
         942 => 8X"20",
         943 => 8X"20",
         944 => 8X"20",
         945 => 8X"20",
         946 => 8X"20",
         947 => 8X"20",
         948 => 8X"20",
         949 => 8X"20",
         950 => 8X"20",
         951 => 8X"20",
         952 => 8X"20",
         953 => 8X"20",
         954 => 8X"20",
         955 => 8X"20",
         956 => 8X"20",
         957 => 8X"20",
         958 => 8X"20",
         959 => 8X"20",
         960 => 8X"74",
         961 => 8X"34",
         962 => 8X"3A",
         963 => 8X"20",
         964 => 8X"30",
         965 => 8X"78",
         966 => 8X"2A",
         967 => 8X"2A",
         968 => 8X"2A",
         969 => 8X"2A",
         970 => 8X"2A",
         971 => 8X"2A",
         972 => 8X"2A",
         973 => 8X"2A",
         974 => 8X"20",
         975 => 8X"20",
         976 => 8X"20",
         977 => 8X"20",
         978 => 8X"20",
         979 => 8X"20",
         980 => 8X"20",
         981 => 8X"20",
         982 => 8X"20",
         983 => 8X"20",
         984 => 8X"20",
         985 => 8X"20",
         986 => 8X"20",
         987 => 8X"20",
         988 => 8X"20",
         989 => 8X"20",
         990 => 8X"20",
         991 => 8X"20",
         992 => 8X"20",
         993 => 8X"20",
         994 => 8X"20",
         995 => 8X"20",
         996 => 8X"20",
         997 => 8X"20",
         998 => 8X"20",
         999 => 8X"20",
        1000 => 8X"20",
        1001 => 8X"20",
        1002 => 8X"20",
        1003 => 8X"20",
        1004 => 8X"20",
        1005 => 8X"20",
        1006 => 8X"20",
        1007 => 8X"20",
        1008 => 8X"20",
        1009 => 8X"20",
        1010 => 8X"20",
        1011 => 8X"20",
        1012 => 8X"20",
        1013 => 8X"20",
        1014 => 8X"20",
        1015 => 8X"20",
        1016 => 8X"20",
        1017 => 8X"20",
        1018 => 8X"20",
        1019 => 8X"20",
        1020 => 8X"20",
        1021 => 8X"20",
        1022 => 8X"20",
        1023 => 8X"20",
        1024 => 8X"20",
        1025 => 8X"20",
        1026 => 8X"20",
        1027 => 8X"20",
        1028 => 8X"20",
        1029 => 8X"20",
        1030 => 8X"20",
        1031 => 8X"20",
        1032 => 8X"20",
        1033 => 8X"20",
        1034 => 8X"20",
        1035 => 8X"20",
        1036 => 8X"20",
        1037 => 8X"20",
        1038 => 8X"20",
        1039 => 8X"20",
        1040 => 8X"74",
        1041 => 8X"35",
        1042 => 8X"3A",
        1043 => 8X"20",
        1044 => 8X"30",
        1045 => 8X"78",
        1046 => 8X"2A",
        1047 => 8X"2A",
        1048 => 8X"2A",
        1049 => 8X"2A",
        1050 => 8X"2A",
        1051 => 8X"2A",
        1052 => 8X"2A",
        1053 => 8X"2A",
        1054 => 8X"20",
        1055 => 8X"20",
        1056 => 8X"20",
        1057 => 8X"20",
        1058 => 8X"20",
        1059 => 8X"20",
        1060 => 8X"20",
        1061 => 8X"20",
        1062 => 8X"20",
        1063 => 8X"20",
        1064 => 8X"20",
        1065 => 8X"20",
        1066 => 8X"20",
        1067 => 8X"20",
        1068 => 8X"20",
        1069 => 8X"20",
        1070 => 8X"20",
        1071 => 8X"20",
        1072 => 8X"20",
        1073 => 8X"20",
        1074 => 8X"20",
        1075 => 8X"20",
        1076 => 8X"20",
        1077 => 8X"20",
        1078 => 8X"20",
        1079 => 8X"20",
        1080 => 8X"20",
        1081 => 8X"20",
        1082 => 8X"20",
        1083 => 8X"20",
        1084 => 8X"20",
        1085 => 8X"20",
        1086 => 8X"20",
        1087 => 8X"20",
        1088 => 8X"20",
        1089 => 8X"20",
        1090 => 8X"20",
        1091 => 8X"20",
        1092 => 8X"20",
        1093 => 8X"20",
        1094 => 8X"20",
        1095 => 8X"20",
        1096 => 8X"20",
        1097 => 8X"20",
        1098 => 8X"20",
        1099 => 8X"20",
        1100 => 8X"20",
        1101 => 8X"20",
        1102 => 8X"20",
        1103 => 8X"20",
        1104 => 8X"20",
        1105 => 8X"20",
        1106 => 8X"20",
        1107 => 8X"20",
        1108 => 8X"20",
        1109 => 8X"20",
        1110 => 8X"20",
        1111 => 8X"20",
        1112 => 8X"20",
        1113 => 8X"20",
        1114 => 8X"20",
        1115 => 8X"20",
        1116 => 8X"20",
        1117 => 8X"20",
        1118 => 8X"20",
        1119 => 8X"20",
        1120 => 8X"74",
        1121 => 8X"36",
        1122 => 8X"3A",
        1123 => 8X"20",
        1124 => 8X"30",
        1125 => 8X"78",
        1126 => 8X"2A",
        1127 => 8X"2A",
        1128 => 8X"2A",
        1129 => 8X"2A",
        1130 => 8X"2A",
        1131 => 8X"2A",
        1132 => 8X"2A",
        1133 => 8X"2A",
        1134 => 8X"20",
        1135 => 8X"20",
        1136 => 8X"20",
        1137 => 8X"20",
        1138 => 8X"20",
        1139 => 8X"20",
        1140 => 8X"20",
        1141 => 8X"20",
        1142 => 8X"20",
        1143 => 8X"20",
        1144 => 8X"20",
        1145 => 8X"20",
        1146 => 8X"20",
        1147 => 8X"20",
        1148 => 8X"20",
        1149 => 8X"20",
        1150 => 8X"20",
        1151 => 8X"20",
        1152 => 8X"20",
        1153 => 8X"20",
        1154 => 8X"20",
        1155 => 8X"20",
        1156 => 8X"20",
        1157 => 8X"20",
        1158 => 8X"20",
        1159 => 8X"20",
        1160 => 8X"20",
        1161 => 8X"20",
        1162 => 8X"20",
        1163 => 8X"20",
        1164 => 8X"20",
        1165 => 8X"20",
        1166 => 8X"20",
        1167 => 8X"20",
        1168 => 8X"20",
        1169 => 8X"20",
        1170 => 8X"20",
        1171 => 8X"20",
        1172 => 8X"20",
        1173 => 8X"20",
        1174 => 8X"20",
        1175 => 8X"20",
        1176 => 8X"20",
        1177 => 8X"20",
        1178 => 8X"20",
        1179 => 8X"20",
        1180 => 8X"20",
        1181 => 8X"20",
        1182 => 8X"20",
        1183 => 8X"20",
        1184 => 8X"20",
        1185 => 8X"20",
        1186 => 8X"20",
        1187 => 8X"20",
        1188 => 8X"20",
        1189 => 8X"20",
        1190 => 8X"20",
        1191 => 8X"20",
        1192 => 8X"20",
        1193 => 8X"20",
        1194 => 8X"20",
        1195 => 8X"20",
        1196 => 8X"20",
        1197 => 8X"20",
        1198 => 8X"20",
        1199 => 8X"20",
        1200 => 8X"74",
        1201 => 8X"37",
        1202 => 8X"3A",
        1203 => 8X"20",
        1204 => 8X"30",
        1205 => 8X"78",
        1206 => 8X"2A",
        1207 => 8X"2A",
        1208 => 8X"2A",
        1209 => 8X"2A",
        1210 => 8X"2A",
        1211 => 8X"2A",
        1212 => 8X"2A",
        1213 => 8X"2A",
        1214 => 8X"20",
        1215 => 8X"20",
        1216 => 8X"20",
        1217 => 8X"20",
        1218 => 8X"20",
        1219 => 8X"20",
        1220 => 8X"20",
        1221 => 8X"20",
        1222 => 8X"20",
        1223 => 8X"20",
        1224 => 8X"20",
        1225 => 8X"20",
        1226 => 8X"20",
        1227 => 8X"20",
        1228 => 8X"20",
        1229 => 8X"20",
        1230 => 8X"20",
        1231 => 8X"20",
        1232 => 8X"20",
        1233 => 8X"20",
        1234 => 8X"20",
        1235 => 8X"20",
        1236 => 8X"20",
        1237 => 8X"20",
        1238 => 8X"20",
        1239 => 8X"20",
        1240 => 8X"20",
        1241 => 8X"20",
        1242 => 8X"20",
        1243 => 8X"20",
        1244 => 8X"20",
        1245 => 8X"20",
        1246 => 8X"20",
        1247 => 8X"20",
        1248 => 8X"20",
        1249 => 8X"20",
        1250 => 8X"20",
        1251 => 8X"20",
        1252 => 8X"20",
        1253 => 8X"20",
        1254 => 8X"20",
        1255 => 8X"20",
        1256 => 8X"20",
        1257 => 8X"20",
        1258 => 8X"20",
        1259 => 8X"20",
        1260 => 8X"20",
        1261 => 8X"20",
        1262 => 8X"20",
        1263 => 8X"20",
        1264 => 8X"20",
        1265 => 8X"20",
        1266 => 8X"20",
        1267 => 8X"20",
        1268 => 8X"20",
        1269 => 8X"20",
        1270 => 8X"20",
        1271 => 8X"20",
        1272 => 8X"20",
        1273 => 8X"20",
        1274 => 8X"20",
        1275 => 8X"20",
        1276 => 8X"20",
        1277 => 8X"20",
        1278 => 8X"20",
        1279 => 8X"20",
        1280 => 8X"73",
        1281 => 8X"30",
        1282 => 8X"3A",
        1283 => 8X"20",
        1284 => 8X"30",
        1285 => 8X"78",
        1286 => 8X"2A",
        1287 => 8X"2A",
        1288 => 8X"2A",
        1289 => 8X"2A",
        1290 => 8X"2A",
        1291 => 8X"2A",
        1292 => 8X"2A",
        1293 => 8X"2A",
        1294 => 8X"20",
        1295 => 8X"20",
        1296 => 8X"20",
        1297 => 8X"20",
        1298 => 8X"20",
        1299 => 8X"20",
        1300 => 8X"20",
        1301 => 8X"20",
        1302 => 8X"20",
        1303 => 8X"20",
        1304 => 8X"20",
        1305 => 8X"20",
        1306 => 8X"20",
        1307 => 8X"20",
        1308 => 8X"20",
        1309 => 8X"20",
        1310 => 8X"20",
        1311 => 8X"20",
        1312 => 8X"20",
        1313 => 8X"20",
        1314 => 8X"20",
        1315 => 8X"20",
        1316 => 8X"20",
        1317 => 8X"20",
        1318 => 8X"20",
        1319 => 8X"20",
        1320 => 8X"20",
        1321 => 8X"20",
        1322 => 8X"20",
        1323 => 8X"20",
        1324 => 8X"20",
        1325 => 8X"20",
        1326 => 8X"20",
        1327 => 8X"20",
        1328 => 8X"20",
        1329 => 8X"20",
        1330 => 8X"20",
        1331 => 8X"20",
        1332 => 8X"20",
        1333 => 8X"20",
        1334 => 8X"20",
        1335 => 8X"20",
        1336 => 8X"20",
        1337 => 8X"20",
        1338 => 8X"20",
        1339 => 8X"20",
        1340 => 8X"20",
        1341 => 8X"20",
        1342 => 8X"20",
        1343 => 8X"20",
        1344 => 8X"20",
        1345 => 8X"20",
        1346 => 8X"20",
        1347 => 8X"20",
        1348 => 8X"20",
        1349 => 8X"20",
        1350 => 8X"20",
        1351 => 8X"20",
        1352 => 8X"20",
        1353 => 8X"20",
        1354 => 8X"20",
        1355 => 8X"20",
        1356 => 8X"20",
        1357 => 8X"20",
        1358 => 8X"20",
        1359 => 8X"20",
        1360 => 8X"73",
        1361 => 8X"31",
        1362 => 8X"3A",
        1363 => 8X"20",
        1364 => 8X"30",
        1365 => 8X"78",
        1366 => 8X"2A",
        1367 => 8X"2A",
        1368 => 8X"2A",
        1369 => 8X"2A",
        1370 => 8X"2A",
        1371 => 8X"2A",
        1372 => 8X"2A",
        1373 => 8X"2A",
        1374 => 8X"20",
        1375 => 8X"20",
        1376 => 8X"20",
        1377 => 8X"20",
        1378 => 8X"20",
        1379 => 8X"20",
        1380 => 8X"20",
        1381 => 8X"20",
        1382 => 8X"20",
        1383 => 8X"20",
        1384 => 8X"20",
        1385 => 8X"20",
        1386 => 8X"20",
        1387 => 8X"20",
        1388 => 8X"20",
        1389 => 8X"20",
        1390 => 8X"20",
        1391 => 8X"20",
        1392 => 8X"20",
        1393 => 8X"20",
        1394 => 8X"20",
        1395 => 8X"20",
        1396 => 8X"20",
        1397 => 8X"20",
        1398 => 8X"20",
        1399 => 8X"20",
        1400 => 8X"20",
        1401 => 8X"20",
        1402 => 8X"20",
        1403 => 8X"20",
        1404 => 8X"20",
        1405 => 8X"20",
        1406 => 8X"20",
        1407 => 8X"20",
        1408 => 8X"20",
        1409 => 8X"20",
        1410 => 8X"20",
        1411 => 8X"20",
        1412 => 8X"20",
        1413 => 8X"20",
        1414 => 8X"20",
        1415 => 8X"20",
        1416 => 8X"20",
        1417 => 8X"20",
        1418 => 8X"20",
        1419 => 8X"20",
        1420 => 8X"20",
        1421 => 8X"20",
        1422 => 8X"20",
        1423 => 8X"20",
        1424 => 8X"20",
        1425 => 8X"20",
        1426 => 8X"20",
        1427 => 8X"20",
        1428 => 8X"20",
        1429 => 8X"20",
        1430 => 8X"20",
        1431 => 8X"20",
        1432 => 8X"20",
        1433 => 8X"20",
        1434 => 8X"20",
        1435 => 8X"20",
        1436 => 8X"20",
        1437 => 8X"20",
        1438 => 8X"20",
        1439 => 8X"20",
        1440 => 8X"73",
        1441 => 8X"32",
        1442 => 8X"3A",
        1443 => 8X"20",
        1444 => 8X"30",
        1445 => 8X"78",
        1446 => 8X"2A",
        1447 => 8X"2A",
        1448 => 8X"2A",
        1449 => 8X"2A",
        1450 => 8X"2A",
        1451 => 8X"2A",
        1452 => 8X"2A",
        1453 => 8X"2A",
        1454 => 8X"20",
        1455 => 8X"20",
        1456 => 8X"20",
        1457 => 8X"20",
        1458 => 8X"20",
        1459 => 8X"20",
        1460 => 8X"20",
        1461 => 8X"20",
        1462 => 8X"20",
        1463 => 8X"20",
        1464 => 8X"20",
        1465 => 8X"20",
        1466 => 8X"20",
        1467 => 8X"20",
        1468 => 8X"20",
        1469 => 8X"20",
        1470 => 8X"20",
        1471 => 8X"20",
        1472 => 8X"20",
        1473 => 8X"20",
        1474 => 8X"20",
        1475 => 8X"20",
        1476 => 8X"20",
        1477 => 8X"20",
        1478 => 8X"20",
        1479 => 8X"20",
        1480 => 8X"20",
        1481 => 8X"20",
        1482 => 8X"20",
        1483 => 8X"20",
        1484 => 8X"20",
        1485 => 8X"20",
        1486 => 8X"20",
        1487 => 8X"20",
        1488 => 8X"20",
        1489 => 8X"20",
        1490 => 8X"20",
        1491 => 8X"20",
        1492 => 8X"20",
        1493 => 8X"20",
        1494 => 8X"20",
        1495 => 8X"20",
        1496 => 8X"20",
        1497 => 8X"20",
        1498 => 8X"20",
        1499 => 8X"20",
        1500 => 8X"20",
        1501 => 8X"20",
        1502 => 8X"20",
        1503 => 8X"20",
        1504 => 8X"20",
        1505 => 8X"20",
        1506 => 8X"20",
        1507 => 8X"20",
        1508 => 8X"20",
        1509 => 8X"20",
        1510 => 8X"20",
        1511 => 8X"20",
        1512 => 8X"20",
        1513 => 8X"20",
        1514 => 8X"20",
        1515 => 8X"20",
        1516 => 8X"20",
        1517 => 8X"20",
        1518 => 8X"20",
        1519 => 8X"20",
        1520 => 8X"73",
        1521 => 8X"33",
        1522 => 8X"3A",
        1523 => 8X"20",
        1524 => 8X"30",
        1525 => 8X"78",
        1526 => 8X"2A",
        1527 => 8X"2A",
        1528 => 8X"2A",
        1529 => 8X"2A",
        1530 => 8X"2A",
        1531 => 8X"2A",
        1532 => 8X"2A",
        1533 => 8X"2A",
        1534 => 8X"20",
        1535 => 8X"20",
        1536 => 8X"20",
        1537 => 8X"20",
        1538 => 8X"20",
        1539 => 8X"20",
        1540 => 8X"20",
        1541 => 8X"20",
        1542 => 8X"20",
        1543 => 8X"20",
        1544 => 8X"20",
        1545 => 8X"20",
        1546 => 8X"20",
        1547 => 8X"20",
        1548 => 8X"20",
        1549 => 8X"20",
        1550 => 8X"20",
        1551 => 8X"20",
        1552 => 8X"20",
        1553 => 8X"20",
        1554 => 8X"20",
        1555 => 8X"20",
        1556 => 8X"20",
        1557 => 8X"20",
        1558 => 8X"20",
        1559 => 8X"20",
        1560 => 8X"20",
        1561 => 8X"20",
        1562 => 8X"20",
        1563 => 8X"20",
        1564 => 8X"20",
        1565 => 8X"20",
        1566 => 8X"20",
        1567 => 8X"20",
        1568 => 8X"20",
        1569 => 8X"20",
        1570 => 8X"20",
        1571 => 8X"20",
        1572 => 8X"20",
        1573 => 8X"20",
        1574 => 8X"20",
        1575 => 8X"20",
        1576 => 8X"20",
        1577 => 8X"20",
        1578 => 8X"20",
        1579 => 8X"20",
        1580 => 8X"20",
        1581 => 8X"20",
        1582 => 8X"20",
        1583 => 8X"20",
        1584 => 8X"20",
        1585 => 8X"20",
        1586 => 8X"20",
        1587 => 8X"20",
        1588 => 8X"20",
        1589 => 8X"20",
        1590 => 8X"20",
        1591 => 8X"20",
        1592 => 8X"20",
        1593 => 8X"20",
        1594 => 8X"20",
        1595 => 8X"20",
        1596 => 8X"20",
        1597 => 8X"20",
        1598 => 8X"20",
        1599 => 8X"20",
        1600 => 8X"73",
        1601 => 8X"34",
        1602 => 8X"3A",
        1603 => 8X"20",
        1604 => 8X"30",
        1605 => 8X"78",
        1606 => 8X"2A",
        1607 => 8X"2A",
        1608 => 8X"2A",
        1609 => 8X"2A",
        1610 => 8X"2A",
        1611 => 8X"2A",
        1612 => 8X"2A",
        1613 => 8X"2A",
        1614 => 8X"20",
        1615 => 8X"20",
        1616 => 8X"20",
        1617 => 8X"20",
        1618 => 8X"20",
        1619 => 8X"20",
        1620 => 8X"20",
        1621 => 8X"20",
        1622 => 8X"20",
        1623 => 8X"20",
        1624 => 8X"20",
        1625 => 8X"20",
        1626 => 8X"20",
        1627 => 8X"20",
        1628 => 8X"20",
        1629 => 8X"20",
        1630 => 8X"20",
        1631 => 8X"20",
        1632 => 8X"20",
        1633 => 8X"20",
        1634 => 8X"20",
        1635 => 8X"20",
        1636 => 8X"20",
        1637 => 8X"20",
        1638 => 8X"20",
        1639 => 8X"20",
        1640 => 8X"20",
        1641 => 8X"20",
        1642 => 8X"20",
        1643 => 8X"20",
        1644 => 8X"20",
        1645 => 8X"20",
        1646 => 8X"20",
        1647 => 8X"20",
        1648 => 8X"20",
        1649 => 8X"20",
        1650 => 8X"20",
        1651 => 8X"20",
        1652 => 8X"20",
        1653 => 8X"20",
        1654 => 8X"20",
        1655 => 8X"20",
        1656 => 8X"20",
        1657 => 8X"20",
        1658 => 8X"20",
        1659 => 8X"20",
        1660 => 8X"20",
        1661 => 8X"20",
        1662 => 8X"20",
        1663 => 8X"20",
        1664 => 8X"20",
        1665 => 8X"20",
        1666 => 8X"20",
        1667 => 8X"20",
        1668 => 8X"20",
        1669 => 8X"20",
        1670 => 8X"20",
        1671 => 8X"20",
        1672 => 8X"20",
        1673 => 8X"20",
        1674 => 8X"20",
        1675 => 8X"20",
        1676 => 8X"20",
        1677 => 8X"20",
        1678 => 8X"20",
        1679 => 8X"20",
        1680 => 8X"73",
        1681 => 8X"35",
        1682 => 8X"3A",
        1683 => 8X"20",
        1684 => 8X"30",
        1685 => 8X"78",
        1686 => 8X"2A",
        1687 => 8X"2A",
        1688 => 8X"2A",
        1689 => 8X"2A",
        1690 => 8X"2A",
        1691 => 8X"2A",
        1692 => 8X"2A",
        1693 => 8X"2A",
        1694 => 8X"20",
        1695 => 8X"20",
        1696 => 8X"20",
        1697 => 8X"20",
        1698 => 8X"20",
        1699 => 8X"20",
        1700 => 8X"20",
        1701 => 8X"20",
        1702 => 8X"20",
        1703 => 8X"20",
        1704 => 8X"20",
        1705 => 8X"20",
        1706 => 8X"20",
        1707 => 8X"20",
        1708 => 8X"20",
        1709 => 8X"20",
        1710 => 8X"20",
        1711 => 8X"20",
        1712 => 8X"20",
        1713 => 8X"20",
        1714 => 8X"20",
        1715 => 8X"20",
        1716 => 8X"20",
        1717 => 8X"20",
        1718 => 8X"20",
        1719 => 8X"20",
        1720 => 8X"20",
        1721 => 8X"20",
        1722 => 8X"20",
        1723 => 8X"20",
        1724 => 8X"20",
        1725 => 8X"20",
        1726 => 8X"20",
        1727 => 8X"20",
        1728 => 8X"20",
        1729 => 8X"20",
        1730 => 8X"20",
        1731 => 8X"20",
        1732 => 8X"20",
        1733 => 8X"20",
        1734 => 8X"20",
        1735 => 8X"20",
        1736 => 8X"20",
        1737 => 8X"20",
        1738 => 8X"20",
        1739 => 8X"20",
        1740 => 8X"20",
        1741 => 8X"20",
        1742 => 8X"20",
        1743 => 8X"20",
        1744 => 8X"20",
        1745 => 8X"20",
        1746 => 8X"20",
        1747 => 8X"20",
        1748 => 8X"20",
        1749 => 8X"20",
        1750 => 8X"20",
        1751 => 8X"20",
        1752 => 8X"20",
        1753 => 8X"20",
        1754 => 8X"20",
        1755 => 8X"20",
        1756 => 8X"20",
        1757 => 8X"20",
        1758 => 8X"20",
        1759 => 8X"20",
        1760 => 8X"73",
        1761 => 8X"36",
        1762 => 8X"3A",
        1763 => 8X"20",
        1764 => 8X"30",
        1765 => 8X"78",
        1766 => 8X"2A",
        1767 => 8X"2A",
        1768 => 8X"2A",
        1769 => 8X"2A",
        1770 => 8X"2A",
        1771 => 8X"2A",
        1772 => 8X"2A",
        1773 => 8X"2A",
        1774 => 8X"20",
        1775 => 8X"20",
        1776 => 8X"20",
        1777 => 8X"20",
        1778 => 8X"20",
        1779 => 8X"20",
        1780 => 8X"20",
        1781 => 8X"20",
        1782 => 8X"20",
        1783 => 8X"20",
        1784 => 8X"20",
        1785 => 8X"20",
        1786 => 8X"20",
        1787 => 8X"20",
        1788 => 8X"20",
        1789 => 8X"20",
        1790 => 8X"20",
        1791 => 8X"20",
        1792 => 8X"20",
        1793 => 8X"20",
        1794 => 8X"20",
        1795 => 8X"20",
        1796 => 8X"20",
        1797 => 8X"20",
        1798 => 8X"20",
        1799 => 8X"20",
        1800 => 8X"20",
        1801 => 8X"20",
        1802 => 8X"20",
        1803 => 8X"20",
        1804 => 8X"20",
        1805 => 8X"20",
        1806 => 8X"20",
        1807 => 8X"20",
        1808 => 8X"20",
        1809 => 8X"20",
        1810 => 8X"20",
        1811 => 8X"20",
        1812 => 8X"20",
        1813 => 8X"20",
        1814 => 8X"20",
        1815 => 8X"20",
        1816 => 8X"20",
        1817 => 8X"20",
        1818 => 8X"20",
        1819 => 8X"20",
        1820 => 8X"20",
        1821 => 8X"20",
        1822 => 8X"20",
        1823 => 8X"20",
        1824 => 8X"20",
        1825 => 8X"20",
        1826 => 8X"20",
        1827 => 8X"20",
        1828 => 8X"20",
        1829 => 8X"20",
        1830 => 8X"20",
        1831 => 8X"20",
        1832 => 8X"20",
        1833 => 8X"20",
        1834 => 8X"20",
        1835 => 8X"20",
        1836 => 8X"20",
        1837 => 8X"20",
        1838 => 8X"20",
        1839 => 8X"20",
        1840 => 8X"73",
        1841 => 8X"37",
        1842 => 8X"3A",
        1843 => 8X"20",
        1844 => 8X"30",
        1845 => 8X"78",
        1846 => 8X"2A",
        1847 => 8X"2A",
        1848 => 8X"2A",
        1849 => 8X"2A",
        1850 => 8X"2A",
        1851 => 8X"2A",
        1852 => 8X"2A",
        1853 => 8X"2A",
        1854 => 8X"20",
        1855 => 8X"20",
        1856 => 8X"20",
        1857 => 8X"20",
        1858 => 8X"20",
        1859 => 8X"20",
        1860 => 8X"20",
        1861 => 8X"20",
        1862 => 8X"20",
        1863 => 8X"20",
        1864 => 8X"20",
        1865 => 8X"20",
        1866 => 8X"20",
        1867 => 8X"20",
        1868 => 8X"20",
        1869 => 8X"20",
        1870 => 8X"20",
        1871 => 8X"20",
        1872 => 8X"20",
        1873 => 8X"20",
        1874 => 8X"20",
        1875 => 8X"20",
        1876 => 8X"20",
        1877 => 8X"20",
        1878 => 8X"20",
        1879 => 8X"20",
        1880 => 8X"20",
        1881 => 8X"20",
        1882 => 8X"20",
        1883 => 8X"20",
        1884 => 8X"20",
        1885 => 8X"20",
        1886 => 8X"20",
        1887 => 8X"20",
        1888 => 8X"20",
        1889 => 8X"20",
        1890 => 8X"20",
        1891 => 8X"20",
        1892 => 8X"20",
        1893 => 8X"20",
        1894 => 8X"20",
        1895 => 8X"20",
        1896 => 8X"20",
        1897 => 8X"20",
        1898 => 8X"20",
        1899 => 8X"20",
        1900 => 8X"20",
        1901 => 8X"20",
        1902 => 8X"20",
        1903 => 8X"20",
        1904 => 8X"20",
        1905 => 8X"20",
        1906 => 8X"20",
        1907 => 8X"20",
        1908 => 8X"20",
        1909 => 8X"20",
        1910 => 8X"20",
        1911 => 8X"20",
        1912 => 8X"20",
        1913 => 8X"20",
        1914 => 8X"20",
        1915 => 8X"20",
        1916 => 8X"20",
        1917 => 8X"20",
        1918 => 8X"20",
        1919 => 8X"20",
        1920 => 8X"74",
        1921 => 8X"38",
        1922 => 8X"3A",
        1923 => 8X"20",
        1924 => 8X"30",
        1925 => 8X"78",
        1926 => 8X"2A",
        1927 => 8X"2A",
        1928 => 8X"2A",
        1929 => 8X"2A",
        1930 => 8X"2A",
        1931 => 8X"2A",
        1932 => 8X"2A",
        1933 => 8X"2A",
        1934 => 8X"20",
        1935 => 8X"20",
        1936 => 8X"20",
        1937 => 8X"20",
        1938 => 8X"20",
        1939 => 8X"20",
        1940 => 8X"20",
        1941 => 8X"20",
        1942 => 8X"20",
        1943 => 8X"20",
        1944 => 8X"20",
        1945 => 8X"20",
        1946 => 8X"20",
        1947 => 8X"20",
        1948 => 8X"20",
        1949 => 8X"20",
        1950 => 8X"20",
        1951 => 8X"20",
        1952 => 8X"20",
        1953 => 8X"20",
        1954 => 8X"20",
        1955 => 8X"20",
        1956 => 8X"20",
        1957 => 8X"20",
        1958 => 8X"20",
        1959 => 8X"20",
        1960 => 8X"20",
        1961 => 8X"20",
        1962 => 8X"20",
        1963 => 8X"20",
        1964 => 8X"20",
        1965 => 8X"20",
        1966 => 8X"20",
        1967 => 8X"20",
        1968 => 8X"20",
        1969 => 8X"20",
        1970 => 8X"20",
        1971 => 8X"20",
        1972 => 8X"20",
        1973 => 8X"20",
        1974 => 8X"20",
        1975 => 8X"20",
        1976 => 8X"20",
        1977 => 8X"20",
        1978 => 8X"20",
        1979 => 8X"20",
        1980 => 8X"20",
        1981 => 8X"20",
        1982 => 8X"20",
        1983 => 8X"20",
        1984 => 8X"20",
        1985 => 8X"20",
        1986 => 8X"20",
        1987 => 8X"20",
        1988 => 8X"20",
        1989 => 8X"20",
        1990 => 8X"20",
        1991 => 8X"20",
        1992 => 8X"20",
        1993 => 8X"20",
        1994 => 8X"20",
        1995 => 8X"20",
        1996 => 8X"20",
        1997 => 8X"20",
        1998 => 8X"20",
        1999 => 8X"20",
        2000 => 8X"74",
        2001 => 8X"39",
        2002 => 8X"3A",
        2003 => 8X"20",
        2004 => 8X"30",
        2005 => 8X"78",
        2006 => 8X"2A",
        2007 => 8X"2A",
        2008 => 8X"2A",
        2009 => 8X"2A",
        2010 => 8X"2A",
        2011 => 8X"2A",
        2012 => 8X"2A",
        2013 => 8X"2A",
        2014 => 8X"20",
        2015 => 8X"20",
        2016 => 8X"20",
        2017 => 8X"20",
        2018 => 8X"20",
        2019 => 8X"20",
        2020 => 8X"20",
        2021 => 8X"20",
        2022 => 8X"20",
        2023 => 8X"20",
        2024 => 8X"20",
        2025 => 8X"20",
        2026 => 8X"20",
        2027 => 8X"20",
        2028 => 8X"20",
        2029 => 8X"20",
        2030 => 8X"20",
        2031 => 8X"20",
        2032 => 8X"20",
        2033 => 8X"20",
        2034 => 8X"20",
        2035 => 8X"20",
        2036 => 8X"20",
        2037 => 8X"20",
        2038 => 8X"20",
        2039 => 8X"20",
        2040 => 8X"20",
        2041 => 8X"20",
        2042 => 8X"20",
        2043 => 8X"20",
        2044 => 8X"20",
        2045 => 8X"20",
        2046 => 8X"20",
        2047 => 8X"20",
        2048 => 8X"20",
        2049 => 8X"20",
        2050 => 8X"20",
        2051 => 8X"20",
        2052 => 8X"20",
        2053 => 8X"20",
        2054 => 8X"20",
        2055 => 8X"20",
        2056 => 8X"20",
        2057 => 8X"20",
        2058 => 8X"20",
        2059 => 8X"20",
        2060 => 8X"20",
        2061 => 8X"20",
        2062 => 8X"20",
        2063 => 8X"20",
        2064 => 8X"20",
        2065 => 8X"20",
        2066 => 8X"20",
        2067 => 8X"20",
        2068 => 8X"20",
        2069 => 8X"20",
        2070 => 8X"20",
        2071 => 8X"20",
        2072 => 8X"20",
        2073 => 8X"20",
        2074 => 8X"20",
        2075 => 8X"20",
        2076 => 8X"20",
        2077 => 8X"20",
        2078 => 8X"20",
        2079 => 8X"20",
        2080 => 8X"6B",
        2081 => 8X"30",
        2082 => 8X"3A",
        2083 => 8X"20",
        2084 => 8X"30",
        2085 => 8X"78",
        2086 => 8X"2A",
        2087 => 8X"2A",
        2088 => 8X"2A",
        2089 => 8X"2A",
        2090 => 8X"2A",
        2091 => 8X"2A",
        2092 => 8X"2A",
        2093 => 8X"2A",
        2094 => 8X"20",
        2095 => 8X"20",
        2096 => 8X"20",
        2097 => 8X"20",
        2098 => 8X"20",
        2099 => 8X"20",
        2100 => 8X"20",
        2101 => 8X"20",
        2102 => 8X"20",
        2103 => 8X"20",
        2104 => 8X"20",
        2105 => 8X"20",
        2106 => 8X"20",
        2107 => 8X"20",
        2108 => 8X"20",
        2109 => 8X"20",
        2110 => 8X"20",
        2111 => 8X"20",
        2112 => 8X"20",
        2113 => 8X"20",
        2114 => 8X"20",
        2115 => 8X"20",
        2116 => 8X"20",
        2117 => 8X"20",
        2118 => 8X"20",
        2119 => 8X"20",
        2120 => 8X"20",
        2121 => 8X"20",
        2122 => 8X"20",
        2123 => 8X"20",
        2124 => 8X"20",
        2125 => 8X"20",
        2126 => 8X"20",
        2127 => 8X"20",
        2128 => 8X"20",
        2129 => 8X"20",
        2130 => 8X"20",
        2131 => 8X"20",
        2132 => 8X"20",
        2133 => 8X"20",
        2134 => 8X"20",
        2135 => 8X"20",
        2136 => 8X"20",
        2137 => 8X"20",
        2138 => 8X"20",
        2139 => 8X"20",
        2140 => 8X"20",
        2141 => 8X"20",
        2142 => 8X"20",
        2143 => 8X"20",
        2144 => 8X"20",
        2145 => 8X"20",
        2146 => 8X"20",
        2147 => 8X"20",
        2148 => 8X"20",
        2149 => 8X"20",
        2150 => 8X"20",
        2151 => 8X"20",
        2152 => 8X"20",
        2153 => 8X"20",
        2154 => 8X"20",
        2155 => 8X"20",
        2156 => 8X"20",
        2157 => 8X"20",
        2158 => 8X"20",
        2159 => 8X"20",
        2160 => 8X"6B",
        2161 => 8X"31",
        2162 => 8X"3A",
        2163 => 8X"20",
        2164 => 8X"30",
        2165 => 8X"78",
        2166 => 8X"2A",
        2167 => 8X"2A",
        2168 => 8X"2A",
        2169 => 8X"2A",
        2170 => 8X"2A",
        2171 => 8X"2A",
        2172 => 8X"2A",
        2173 => 8X"2A",
        2174 => 8X"20",
        2175 => 8X"20",
        2176 => 8X"20",
        2177 => 8X"20",
        2178 => 8X"20",
        2179 => 8X"20",
        2180 => 8X"20",
        2181 => 8X"20",
        2182 => 8X"20",
        2183 => 8X"20",
        2184 => 8X"20",
        2185 => 8X"20",
        2186 => 8X"20",
        2187 => 8X"20",
        2188 => 8X"20",
        2189 => 8X"20",
        2190 => 8X"20",
        2191 => 8X"20",
        2192 => 8X"20",
        2193 => 8X"20",
        2194 => 8X"20",
        2195 => 8X"20",
        2196 => 8X"20",
        2197 => 8X"20",
        2198 => 8X"20",
        2199 => 8X"20",
        2200 => 8X"20",
        2201 => 8X"20",
        2202 => 8X"20",
        2203 => 8X"20",
        2204 => 8X"20",
        2205 => 8X"20",
        2206 => 8X"20",
        2207 => 8X"20",
        2208 => 8X"20",
        2209 => 8X"20",
        2210 => 8X"20",
        2211 => 8X"20",
        2212 => 8X"20",
        2213 => 8X"20",
        2214 => 8X"20",
        2215 => 8X"20",
        2216 => 8X"20",
        2217 => 8X"20",
        2218 => 8X"20",
        2219 => 8X"20",
        2220 => 8X"20",
        2221 => 8X"20",
        2222 => 8X"20",
        2223 => 8X"20",
        2224 => 8X"20",
        2225 => 8X"20",
        2226 => 8X"20",
        2227 => 8X"20",
        2228 => 8X"20",
        2229 => 8X"20",
        2230 => 8X"20",
        2231 => 8X"20",
        2232 => 8X"20",
        2233 => 8X"20",
        2234 => 8X"20",
        2235 => 8X"20",
        2236 => 8X"20",
        2237 => 8X"20",
        2238 => 8X"20",
        2239 => 8X"20",
        2240 => 8X"67",
        2241 => 8X"70",
        2242 => 8X"3A",
        2243 => 8X"20",
        2244 => 8X"30",
        2245 => 8X"78",
        2246 => 8X"2A",
        2247 => 8X"2A",
        2248 => 8X"2A",
        2249 => 8X"2A",
        2250 => 8X"2A",
        2251 => 8X"2A",
        2252 => 8X"2A",
        2253 => 8X"2A",
        2254 => 8X"20",
        2255 => 8X"20",
        2256 => 8X"20",
        2257 => 8X"20",
        2258 => 8X"20",
        2259 => 8X"20",
        2260 => 8X"20",
        2261 => 8X"20",
        2262 => 8X"20",
        2263 => 8X"20",
        2264 => 8X"20",
        2265 => 8X"20",
        2266 => 8X"20",
        2267 => 8X"20",
        2268 => 8X"20",
        2269 => 8X"20",
        2270 => 8X"20",
        2271 => 8X"20",
        2272 => 8X"20",
        2273 => 8X"20",
        2274 => 8X"20",
        2275 => 8X"20",
        2276 => 8X"20",
        2277 => 8X"20",
        2278 => 8X"20",
        2279 => 8X"20",
        2280 => 8X"20",
        2281 => 8X"20",
        2282 => 8X"20",
        2283 => 8X"20",
        2284 => 8X"20",
        2285 => 8X"20",
        2286 => 8X"20",
        2287 => 8X"20",
        2288 => 8X"20",
        2289 => 8X"20",
        2290 => 8X"20",
        2291 => 8X"20",
        2292 => 8X"20",
        2293 => 8X"20",
        2294 => 8X"20",
        2295 => 8X"20",
        2296 => 8X"20",
        2297 => 8X"20",
        2298 => 8X"20",
        2299 => 8X"20",
        2300 => 8X"20",
        2301 => 8X"20",
        2302 => 8X"20",
        2303 => 8X"20",
        2304 => 8X"20",
        2305 => 8X"20",
        2306 => 8X"20",
        2307 => 8X"20",
        2308 => 8X"20",
        2309 => 8X"20",
        2310 => 8X"20",
        2311 => 8X"20",
        2312 => 8X"20",
        2313 => 8X"20",
        2314 => 8X"20",
        2315 => 8X"20",
        2316 => 8X"20",
        2317 => 8X"20",
        2318 => 8X"20",
        2319 => 8X"20",
        2320 => 8X"73",
        2321 => 8X"70",
        2322 => 8X"3A",
        2323 => 8X"20",
        2324 => 8X"30",
        2325 => 8X"78",
        2326 => 8X"2A",
        2327 => 8X"2A",
        2328 => 8X"2A",
        2329 => 8X"2A",
        2330 => 8X"2A",
        2331 => 8X"2A",
        2332 => 8X"2A",
        2333 => 8X"2A",
        2334 => 8X"20",
        2335 => 8X"20",
        2336 => 8X"20",
        2337 => 8X"20",
        2338 => 8X"20",
        2339 => 8X"20",
        2340 => 8X"20",
        2341 => 8X"20",
        2342 => 8X"20",
        2343 => 8X"20",
        2344 => 8X"20",
        2345 => 8X"20",
        2346 => 8X"20",
        2347 => 8X"20",
        2348 => 8X"20",
        2349 => 8X"20",
        2350 => 8X"20",
        2351 => 8X"20",
        2352 => 8X"20",
        2353 => 8X"20",
        2354 => 8X"20",
        2355 => 8X"20",
        2356 => 8X"20",
        2357 => 8X"20",
        2358 => 8X"20",
        2359 => 8X"20",
        2360 => 8X"20",
        2361 => 8X"20",
        2362 => 8X"20",
        2363 => 8X"20",
        2364 => 8X"20",
        2365 => 8X"20",
        2366 => 8X"20",
        2367 => 8X"20",
        2368 => 8X"20",
        2369 => 8X"20",
        2370 => 8X"20",
        2371 => 8X"20",
        2372 => 8X"20",
        2373 => 8X"20",
        2374 => 8X"20",
        2375 => 8X"20",
        2376 => 8X"20",
        2377 => 8X"20",
        2378 => 8X"20",
        2379 => 8X"20",
        2380 => 8X"20",
        2381 => 8X"20",
        2382 => 8X"20",
        2383 => 8X"20",
        2384 => 8X"20",
        2385 => 8X"20",
        2386 => 8X"20",
        2387 => 8X"20",
        2388 => 8X"20",
        2389 => 8X"20",
        2390 => 8X"20",
        2391 => 8X"20",
        2392 => 8X"20",
        2393 => 8X"20",
        2394 => 8X"20",
        2395 => 8X"20",
        2396 => 8X"20",
        2397 => 8X"20",
        2398 => 8X"20",
        2399 => 8X"20",
        2400 => 8X"66",
        2401 => 8X"70",
        2402 => 8X"3A",
        2403 => 8X"20",
        2404 => 8X"30",
        2405 => 8X"78",
        2406 => 8X"2A",
        2407 => 8X"2A",
        2408 => 8X"2A",
        2409 => 8X"2A",
        2410 => 8X"2A",
        2411 => 8X"2A",
        2412 => 8X"2A",
        2413 => 8X"2A",
        2414 => 8X"20",
        2415 => 8X"20",
        2416 => 8X"20",
        2417 => 8X"20",
        2418 => 8X"20",
        2419 => 8X"20",
        2420 => 8X"20",
        2421 => 8X"20",
        2422 => 8X"20",
        2423 => 8X"20",
        2424 => 8X"20",
        2425 => 8X"20",
        2426 => 8X"20",
        2427 => 8X"20",
        2428 => 8X"20",
        2429 => 8X"20",
        2430 => 8X"20",
        2431 => 8X"20",
        2432 => 8X"20",
        2433 => 8X"20",
        2434 => 8X"20",
        2435 => 8X"20",
        2436 => 8X"20",
        2437 => 8X"20",
        2438 => 8X"20",
        2439 => 8X"20",
        2440 => 8X"20",
        2441 => 8X"20",
        2442 => 8X"20",
        2443 => 8X"20",
        2444 => 8X"20",
        2445 => 8X"20",
        2446 => 8X"20",
        2447 => 8X"20",
        2448 => 8X"20",
        2449 => 8X"20",
        2450 => 8X"20",
        2451 => 8X"20",
        2452 => 8X"20",
        2453 => 8X"20",
        2454 => 8X"20",
        2455 => 8X"20",
        2456 => 8X"20",
        2457 => 8X"20",
        2458 => 8X"20",
        2459 => 8X"20",
        2460 => 8X"20",
        2461 => 8X"20",
        2462 => 8X"20",
        2463 => 8X"20",
        2464 => 8X"20",
        2465 => 8X"20",
        2466 => 8X"20",
        2467 => 8X"20",
        2468 => 8X"20",
        2469 => 8X"20",
        2470 => 8X"20",
        2471 => 8X"20",
        2472 => 8X"20",
        2473 => 8X"20",
        2474 => 8X"20",
        2475 => 8X"20",
        2476 => 8X"20",
        2477 => 8X"20",
        2478 => 8X"20",
        2479 => 8X"20",
        2480 => 8X"72",
        2481 => 8X"61",
        2482 => 8X"3A",
        2483 => 8X"20",
        2484 => 8X"30",
        2485 => 8X"78",
        2486 => 8X"2A",
        2487 => 8X"2A",
        2488 => 8X"2A",
        2489 => 8X"2A",
        2490 => 8X"2A",
        2491 => 8X"2A",
        2492 => 8X"2A",
        2493 => 8X"2A",
        2494 => 8X"20",
        2495 => 8X"20",
        2496 => 8X"20",
        2497 => 8X"20",
        2498 => 8X"20",
        2499 => 8X"20",
        2500 => 8X"20",
        2501 => 8X"20",
        2502 => 8X"20",
        2503 => 8X"20",
        2504 => 8X"20",
        2505 => 8X"20",
        2506 => 8X"20",
        2507 => 8X"20",
        2508 => 8X"20",
        2509 => 8X"20",
        2510 => 8X"20",
        2511 => 8X"20",
        2512 => 8X"20",
        2513 => 8X"20",
        2514 => 8X"20",
        2515 => 8X"20",
        2516 => 8X"20",
        2517 => 8X"20",
        2518 => 8X"20",
        2519 => 8X"20",
        2520 => 8X"20",
        2521 => 8X"20",
        2522 => 8X"20",
        2523 => 8X"20",
        2524 => 8X"20",
        2525 => 8X"20",
        2526 => 8X"20",
        2527 => 8X"20",
        2528 => 8X"20",
        2529 => 8X"20",
        2530 => 8X"20",
        2531 => 8X"20",
        2532 => 8X"20",
        2533 => 8X"20",
        2534 => 8X"20",
        2535 => 8X"20",
        2536 => 8X"20",
        2537 => 8X"20",
        2538 => 8X"20",
        2539 => 8X"20",
        2540 => 8X"20",
        2541 => 8X"20",
        2542 => 8X"20",
        2543 => 8X"20",
        2544 => 8X"20",
        2545 => 8X"20",
        2546 => 8X"20",
        2547 => 8X"20",
        2548 => 8X"20",
        2549 => 8X"20",
        2550 => 8X"20",
        2551 => 8X"20",
        2552 => 8X"20",
        2553 => 8X"20",
        2554 => 8X"20",
        2555 => 8X"20",
        2556 => 8X"20",
        2557 => 8X"20",
        2558 => 8X"20",
        2559 => 8X"20",
        others => X"XX"
    );

end package display_mem_schoolMIPS_pkg;
